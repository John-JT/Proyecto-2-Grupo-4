`timescale 1ns / 1ps

// ROM with synchonous read (inferring Block RAM)
// character ROM
//  - 8-by-16 (8-by-2^4) font
//  - 128 (2^7) characters
//  - ROM size: 512-by-8 (2^11-by-8) bits
//              16K bits: 1 BRAM

module font_rom8x16
   (
    input wire [9:0] Qh,
    input wire [9:0] Qv,
    input wire resetM,
    input wire reloj,
    output wire BIT_FUENTE2
   );
   
   // signal declaration
   reg [19:0] addr_reg;
   reg [15:0] data; 
   wire[19:0] addr;
   reg [3:0] SELEC_PX;
   reg bit_fuente2;
   
   Posicion_ROM8x16 inst_Posicion_ROM8x16(
   .resetM(resetM),
   .Qh(Qh[9:3]),
   .Qv(Qv),
   .reloj(reloj),
   .DIR8x16 (addr)
   );

   // body
    always @(*) begin
      SELEC_PX <= {Qh[3], Qh[2], Qh[1], Qh[0]};
      end
   always @(posedge reloj) 
      addr_reg <= addr;
      
   always @*
      case (addr_reg)
         //code x000
         20'h00000: data = 16'h0000; // 
         20'h00001: data = 16'h0000; // 
         20'h00002: data = 16'h0000; // 
         20'h00003: data = 16'h0000; // 
         20'h00004: data = 16'h0000; // 
         20'h00005: data = 16'h0000; // 
         20'h00006: data = 16'h0000; // 
         20'h00007: data = 16'h0000; // 
         20'h00008: data = 16'h0000; // 
         20'h00009: data = 16'h0000; // 
         20'h0000a: data = 16'h0000; // 
         20'h0000b: data = 16'h0000; // 
         20'h0000c: data = 16'h0000; // 
         20'h0000d: data = 16'h0000; // 
         20'h0000e: data = 16'h0000; // 
         20'h0000f: data = 16'h0000; // 
         20'h00010: data = 16'h0000; // 
         20'h00011: data = 16'h0000; // 
         20'h00012: data = 16'h0000; //
         20'h00013: data = 16'h0000; //
         20'h00014: data = 16'h0000; //
         20'h00015: data = 16'h0000; //
         20'h00016: data = 16'h0000; //
         20'h00017: data = 16'h0000; //
         20'h00018: data = 16'h0000; //
         20'h00019: data = 16'h0000; //
         20'h0001a: data = 16'h0000; //
         20'h0001b: data = 16'h0000; //
         20'h0001c: data = 16'h0000; //
         20'h0001d: data = 16'h0000; // 
         20'h0001e: data = 16'h0000; // 
         20'h0001f: data = 16'h0000; // 
         
         /*0*/
         //code x010
         20'h01020: data = 	16'h0000; //
         20'h01021: data = 	16'h0000; //               
         20'h01022: data = 	16'h0000; //               
         20'h01023: data = 	16'h0000; //               
         20'h01024: data = 	16'h0000; //                
         20'h01025: data = 	16'h0000; //                
         20'h01026: data = 	16'h0000; //                
         20'h01027: data = 	16'h0000; //                
         20'h01028: data =  16'h00F8; //         *****  
         20'h01029: data = 	16'h03FC; //       ******** 
         20'h0102a: data = 	16'h071C; //      ***   *** 
         20'h0102b: data = 	16'h0C0E; //     **      ***
         20'h0102c: data = 	16'h180E; //    **       ***
         20'h0102d: data = 	16'h300C; //   **        ** 
         20'h0102e: data = 	16'h600C; //  **         ** 
         20'h0102f: data = 	16'h600C; //  **         ** 
         20'h01030: data = 	16'h6008; //  **         *  
         20'h01031: data = 	16'hC018; // **         **  
         20'h01032: data = 	16'hC030; // **        **   
         20'h01033: data = 	16'hC030; // **        **   
         20'h01034: data = 	16'hC060; // **       **    
         20'h01035: data = 	16'hE1C0; // ***    ***     
         20'h01036: data = 	16'h7F80; //  ********      
         20'h01037: data = 	16'h3E00; //   *****        
         20'h01038: data = 	16'h0000; //                
         20'h01039: data = 	16'h0000; //                
         20'h0103a: data = 	16'h0000; //                
         20'h0103b: data = 	16'h0000; //                
         20'h0103c: data = 	16'h0000; // 
         20'h0103d: data = 	16'h0000; //               
         20'h0103e: data = 	16'h0000; //               
         20'h0103f: data = 	16'h0000; //
                        
         /*1*/
         //code x020
         20'h02040: data =	16'h0000; //
         20'h02041: data =	16'h0000; //               
         20'h02042: data =	16'h0000; //               
         20'h02043: data =	16'h0000; //               
         20'h02044: data =	16'h0000; //               
         20'h02045: data =	16'h0000; //            
         20'h02046: data =	16'h0000; //            
         20'h02047: data =	16'h0000; //            
         20'h02048: data =	16'h0000; //            
         20'h02049: data =	16'h00E0; //         ***
         20'h0204a: data =	16'h07E0; //      ******
         20'h0204b: data =	16'h0F60; //     **** **
         20'h0204c: data =	16'h1CC0; //    ***  ** 
         20'h0204d: data =	16'h00C0; //         ** 
         20'h0204e: data =	16'h0180; //        **  
         20'h0204f: data =	16'h0180; //        **  
         20'h02050: data =	16'h0300; //       **   
         20'h02051: data =	16'h0300; //       **   
         20'h02052: data =	16'h0600; //      **    
         20'h02053: data =	16'h0600; //      **    
         20'h02054: data =	16'h0C00; //     **     
         20'h02055: data =	16'h0C00; //     **     
         20'h02056: data =	16'hD800; // ** **      
         20'h02057: data =	16'hFF00; // ********   
         20'h02058: data =	16'h7F00; //  *******   
         20'h02059: data =	16'h0000; //            
         20'h0205a: data =	16'h0000; //            
         20'h0205b: data =	16'h0000; //            
         20'h0205c: data =	16'h0000; //            
         20'h0205d: data =	16'h0000; //
         20'h0205e: data =	16'h0000; //               
         20'h0205f: data =	16'h0000; // 
             
         /*2*/
         //code x030      	              
         20'h03060: data =  16'h0000; //               
         20'h03061: data = 	16'h0000; //               
         20'h03062: data = 	16'h0000; //               
         20'h03063: data = 	16'h0000; //              
         20'h03064: data = 	16'h0000; //              
         20'h03065: data = 	16'h0000; //              
         20'h03066: data = 	16'h0000; //              
         20'h03067: data = 	16'h00F8; //         *****
         20'h03068: data = 	16'h03F8; //       *******
         20'h03069: data = 	16'h0798; //      ****  **
         20'h0306a: data = 	16'h0E18; //     ***    **
         20'h0306b: data = 	16'h0018; //            **
         20'h0306c: data = 	16'h0018; //            **
         20'h0306d: data = 	16'h0030; //           ** 
         20'h0306e: data = 	16'h0060; //          **  
         20'h0306f: data = 	16'h00E0; //         ***  
         20'h03070: data = 	16'h01C0; //        ***   
         20'h03071: data = 	16'h0380; //       ***    
         20'h03072: data = 	16'h0E00; //     ***      
         20'h03073: data = 	16'h1C00; //    ***       
         20'h03074: data = 	16'h7070; //  ***     *** 
         20'h03075: data = 	16'hFFE0; // ***********  
         20'h03076: data = 	16'hFF00; // ********     
         20'h03077: data = 	16'h0000; //              
         20'h03078: data = 	16'h0000; //              
         20'h03079: data = 	16'h0000; //              
         20'h0307a: data = 	16'h0000; //              
         20'h0307b: data = 	16'h0000; //     
         20'h0307c: data = 	16'h0000; //               
         20'h0307d: data = 	16'h0000; //               
         20'h0307e: data = 	16'h0000; //               
         20'h0307f: data = 	16'h0000; // 
                       
         /*3*/
         //code x040
         20'h04080: data = 	16'h0000; //               
         20'h04081: data = 	16'h0000; //               
         20'h04082: data = 	16'h0000; //               
         20'h04083: data = 	16'h0000; //             
         20'h04084: data = 	16'h0000; //             
         20'h04085: data = 	16'h0000; //             
         20'h04086: data = 	16'h0000; //             
         20'h04087: data = 	16'h01E0; //        **** 
         20'h04088: data = 	16'h03F0; //       ******
         20'h04089: data = 	16'h0030; //           **
         20'h0408a: data = 	16'h0030; //           **
         20'h0408b: data = 	16'h0030; //           **
         20'h0408c: data = 	16'h0060; //          ** 
         20'h0408d: data = 	16'h07C0; //      *****  
         20'h0408e: data = 	16'h07C0; //      *****  
         20'h0408f: data = 	16'h00E0; //         *** 
         20'h04090: data = 	16'h0060; //          ** 
         20'h04091: data = 	16'h0060; //          ** 
         20'h04092: data = 	16'h0060; //          ** 
         20'h04093: data = 	16'hC0C0; // **      **  
         20'h04094: data = 	16'hC380; // **    ***   
         20'h04095: data = 	16'hFF00; // ********    
         20'h04096: data = 	16'hFC00; // ******      
         20'h04097: data = 	16'h0000; //             
         20'h04098: data = 	16'h0000; //             
         20'h04099: data = 	16'h0000; //             
         20'h0409a: data = 	16'h0000; //             
         20'h0409b: data = 	16'h0000; // 
         20'h0409c: data = 	16'h0000; //               
         20'h0409d: data = 	16'h0000; //               
         20'h0409e: data = 	16'h0000; //               
         20'h0409f: data = 	16'h0000; //    
                    
         /*4*/
         //code x050
         20'h050a0: data =	16'h0000; //               
         20'h050a1: data =	16'h0000; //               
         20'h050a2: data =	16'h0000; //               
         20'h050a3: data =	16'h0000; //             
         20'h050a4: data =	16'h0000; //             
         20'h050a5: data =	16'h0000; //             
         20'h050a6: data =	16'h0000; //             
         20'h050a7: data =	16'h0300; //       **    
         20'h050a8: data =	16'h0730; //      ***  **
         20'h050a9: data =	16'h0C70; //     **   ***
         20'h050aa: data =	16'h18E0; //    **   *** 
         20'h050ab: data =	16'h30C0; //   **    **  
         20'h050ac: data =	16'h61C0; //  **    ***  
         20'h050ad: data =	16'h4180; //  *     **   
         20'h050ae: data =	16'hC300; // **    **    
         20'h050af: data =	16'hE340; // ***   ** *  
         20'h050b0: data =	16'hFFC0; // **********  
         20'h050b1: data =	16'h7F80; //  ********   
         20'h050b2: data =	16'h0C00; //     **      
         20'h050b3: data =	16'h0800; //     *       
         20'h050b4: data =	16'h1800; //    **       
         20'h050b5: data =	16'h1800; //    **       
         20'h050b6: data =	16'h3000; //   **        
         20'h050b7: data =	16'h3000; //   **        
         20'h050b8: data =	16'h0000; //             
         20'h050b9: data =	16'h0000; //             
         20'h050ba: data =	16'h0000; //             
         20'h050bb: data =	16'h0000; //  
         20'h050bc: data =	16'h0000; //               
         20'h050bd: data =	16'h0000; //               
         20'h050be: data =	16'h0000; //               
         20'h050bf: data =	16'h0000; //  
         
         /*5*/                        
         //code x060         
         20'h060c0: data =  16'h0000; //               
         20'h060c1: data =  16'h0000; //               
         20'h060c2: data =  16'h0000; //               
         20'h060c3: data = 	16'h0000; //               
         20'h060c4: data = 	16'h0000; //               
         20'h060c5: data =  16'h0000; //               
         20'h060c6: data =  16'h01F0; //        *****  
         20'h060c7: data =  16'h03FC; //       ********
         20'h060c8: data =  16'h071C; //      ***   ***
         20'h060c9: data =  16'h0600; //      **       
         20'h060ca: data =  16'h0C00; //     **        
         20'h060cb: data =  16'h0FC0; //     ******    
         20'h060cc: data =  16'h0FF0; //     ********  
         20'h060cd: data =  16'h1870; //    **    ***  
         20'h060ce: data =  16'h0030; //           **  
         20'h060cf: data =  16'h0030; //           **  
         20'h060d0: data =  16'h0030; //           **  
         20'h060d1: data =  16'h0030; //           **  
         20'h060d2: data =  16'h0060; //          **   
         20'h060d3: data =  16'hC060; // **       **   
         20'h060d4: data =  16'hC0C0; // **      **    
         20'h060d5: data =  16'hE180; // ***    **     
         20'h060d6: data =  16'hFF00; // ********      
         20'h060d7: data =  16'h7C00; //  *****        
         20'h060d8: data =  16'h0000; //               
         20'h060d9: data =  16'h0000; //               
         20'h060da: data =  16'h0000; //               
         20'h060db: data = 	16'h0000; // 
         20'h060dc: data = 	16'h0000; //               
         20'h060dd: data =  16'h0000; //               
         20'h060de: data =  16'h0000; //               
         20'h060df: data =  16'h0000; //    
         
         /*6*/                         
         //code x070
         20'h070e0: data = 	16'h0000; //               
         20'h070e1: data = 	16'h0000; //               
         20'h070e2: data = 	16'h0000; //               
         20'h070e3: data = 	16'h0000; //               
         20'h070e4: data = 	16'h0000; //               
         20'h070e5: data = 	16'h0000; //               
         20'h070e6: data = 	16'h0078; //          **** 
         20'h070e7: data = 	16'h01FC; //        *******
         20'h070e8: data = 	16'h031C; //       **   ***
         20'h070e9: data = 	16'h0608; //      **     * 
         20'h070ea: data = 	16'h0C00; //     **        
         20'h070eb: data = 	16'h1800; //    **         
         20'h070ec: data = 	16'h1800; //    **         
         20'h070ed: data = 	16'h3000; //   **          
         20'h070ee: data = 	16'h3780; //   ** ****     
         20'h070ef: data = 	16'h3FC0; //   ********    
         20'h070f0: data = 	16'h70E0; //  ***    ***   
         20'h070f1: data = 	16'h60E0; //  **     ***   
         20'h070f2: data = 	16'h60E0; //  **     ***   
         20'h070f3: data = 	16'hC0C0; // **      **    
         20'h070f4: data = 	16'hC0C0; // **      **    
         20'h070f5: data = 	16'h6180; //  **    **     
         20'h070f6: data = 	16'h7F00; //  *******      
         20'h070f7: data = 	16'h3C00; //   ****        
         20'h070f8: data = 	16'h0000; //               
         20'h070f9: data = 	16'h0000; //               
         20'h070fa: data = 	16'h0000; //               
         20'h070fb: data = 	16'h0000; //
         20'h070fc: data = 	16'h0000; //               
         20'h070fd: data = 	16'h0000; //               
         20'h070fe: data = 	16'h0000; //               
         20'h070ff: data = 	16'h0000; //   
                   
         /*7*/            
         //code x081
         20'h08100: data = 	16'h0000; //               
         20'h08101: data = 	16'h0000; //               
         20'h08102: data = 	16'h0000; //               
         20'h08103: data = 	16'h0000; //                 
         20'h08104: data = 	16'h0000; //                 
         20'h08105: data = 	16'h0000; //                 
         20'h08106: data = 	16'h0000; //                 
         20'h08107: data = 	16'h03FE; //       ********* 
         20'h08108: data = 	16'h0FFF; //     ************
         20'h08109: data = 	16'h0C07; //     **       ***
         20'h0810a: data = 	16'h1806; //    **        ** 
         20'h0810b: data = 	16'h000C; //             **  
         20'h0810c: data = 	16'h0018; //            **   
         20'h0810d: data = 	16'h0038; //           ***   
         20'h0810e: data = 	16'h0030; //           **    
         20'h0810f: data = 	16'h0060; //          **     
         20'h08110: data = 	16'h00C0; //         **      
         20'h08111: data = 	16'h0180; //        **       
         20'h08112: data = 	16'h0700; //      ***        
         20'h08113: data = 	16'h0E00; //     ***         
         20'h08114: data = 	16'h1C00; //    ***          
         20'h08115: data = 	16'h3800; //   ***           
         20'h08116: data = 	16'hF000; // ****            
         20'h08117: data = 	16'hC000; // **              
         20'h08118: data = 	16'h0000; //                 
         20'h08119: data = 	16'h0000; //                 
         20'h0811a: data = 	16'h0000; //                 
         20'h0811b: data = 	16'h0000; // 
         20'h0811c: data = 	16'h0000; //               
         20'h0811d: data = 	16'h0000; //               
         20'h0811e: data = 	16'h0000; //               
         20'h0811f: data = 	16'h0000; //   
         
         /*8*/            
         //code x091            
         20'h09120: data = 	16'h0000; //               
         20'h09121: data = 	16'h0000; //               
         20'h09122: data = 	16'h0000; //               
         20'h09123: data = 	16'h0000; //               
         20'h09124: data = 	16'h0000; //               
         20'h09125: data = 	16'h0000; //               
         20'h09126: data = 	16'h0000; //               
         20'h09127: data = 	16'h00F8; //         ***** 
         20'h09128: data = 	16'h03FC; //       ********
         20'h09129: data = 	16'h071C; //      ***   ***
         20'h0912a: data = 	16'h0C0C; //     **      **
         20'h0912b: data = 	16'h0C0C; //     **      **
         20'h0912c: data = 	16'h0C18; //     **     ** 
         20'h0912d: data = 	16'h0C38; //     **    *** 
         20'h0912e: data = 	16'h0FE0; //     *******   
         20'h0912f: data = 	16'h1FE0; //    ********   
         20'h09130: data = 	16'h3070; //   **     ***  
         20'h09131: data = 	16'h6030; //  **       **  
         20'h09132: data = 	16'h6030; //  **       **  
         20'h09133: data = 	16'hC060; // **       **   
         20'h09134: data = 	16'hE0C0; // ***     **    
         20'h09135: data = 	16'h7F80; //  ********     
         20'h09136: data = 	16'h3E00; //   *****       
         20'h09137: data = 	16'h0000; //               
         20'h09138: data = 	16'h0000; //               
         20'h09139: data = 	16'h0000; //               
         20'h0913a: data = 	16'h0000; //               
         20'h0913b: data = 	16'h0000; //
         20'h0913c: data = 	16'h0000; //               
         20'h0913d: data = 	16'h0000; //               
         20'h0913e: data = 	16'h0000; //               
         20'h0913f: data = 	16'h0000; //
            
         /*9*/            
         //code x0a1
         20'h0a140: data = 	16'h0000; //               
         20'h0a141: data = 	16'h0000; //         
         20'h0a142: data = 	16'h0000; //               
         20'h0a143: data = 	16'h0000; //               
         20'h0a144: data = 	16'h0000; //               
         20'h0a145: data = 	16'h0000; //               
         20'h0a146: data = 	16'h01F0; //        *****  
         20'h0a147: data = 	16'h07F8; //      ******** 
         20'h0a148: data = 	16'h0E1C; //     ***    ***
         20'h0a149: data = 	16'h0C0C; //     **      **
         20'h0a14a: data = 	16'h180C; //    **       **
         20'h0a14b: data = 	16'h180C; //    **       **
         20'h0a14c: data = 	16'h3818; //   ***      ** 
         20'h0a14d: data = 	16'h1878; //    **    **** 
         20'h0a14e: data = 	16'h1FF0; //    *********  
         20'h0a14f: data = 	16'h0FB0; //     ***** **  
         20'h0a150: data = 	16'h0060; //          **   
         20'h0a151: data = 	16'h00C0; //         **    
         20'h0a152: data = 	16'h0180; //        **     
         20'h0a153: data = 	16'h0700; //      ***      
         20'h0a154: data = 	16'h1E00; //    ****       
         20'h0a155: data = 	16'h7C00; //  *****        
         20'h0a156: data = 	16'hF000; // ****          
         20'h0a157: data = 	16'hC000; // **            
         20'h0a158: data = 	16'h0000; //               
         20'h0a159: data = 	16'h0000; //               
         20'h0a15a: data = 	16'h0000; //
         20'h0a15b: data = 	16'h0000; //               
         20'h0a15c: data = 	16'h0000; //               
         20'h0a15d: data = 	16'h0000; //
         20'h0a15e: data = 	16'h0000; //  
         20'h0a15f: data = 	16'h0000; //  
                  
         //code x0b1
         /*A*/
         20'h0b160: data =  16'h0000; //               
         20'h0b161: data =  16'h0000; //               
         20'h0b162: data =  16'h0000; //               
         20'h0b163: data =  16'h0000; //               
         20'h0b164: data =  16'h0600; //      11       
         20'h0b165: data =  16'h0600; //      11       
         20'h0b166: data =  16'h0600; //      11       
         20'h0b167: data =  16'h0600; //      11       
         20'h0b168: data =  16'h0600; //      11       
         20'h0b169: data =  16'h0F00; //     1111      
         20'h0b16a: data =  16'h0F00; //     1111      
         20'h0b16b: data =  16'h0F00; //     1111      
         20'h0b16c: data =  16'h0F00; //     1111      
         20'h0b16d: data =  16'h0F00; //     1111      
         20'h0b16e: data =  16'h0F00; //     1111      
         20'h0b16f: data =  16'h1B80; //    11 111     
         20'h0b170: data =  16'h1980; //    11  11     
         20'h0b171: data =  16'h1F80; //    111111     
         20'h0b172: data =  16'h1980; //    11  11     
         20'h0b173: data =  16'h1980; //    11  11     
         20'h0b174: data =  16'h38C0; //   111   11    
         20'h0b175: data =  16'h38C0; //   111   11    
         20'h0b176: data =  16'h38C0; //   111   11    
         20'h0b177: data =  16'h38C0; //   111   11    
         20'h0b178: data =  16'h30C0; //   11    11    
         20'h0b179: data =  16'h71E0; // 1111   11111  
         20'h0b17a: data =  16'h0000; //               
         20'h0b17b: data =  16'h0000; //               
         20'h0b17c: data =  16'h0000; //               
         20'h0b17d: data =  16'h0000; //               
         20'h0b17e: data =  16'h0000; //               
         20'h0b17f: data =  16'h0000; //  
         
         /*B*/             
         //code x0c1
         20'h0c180: data = 	16'h0000; //               
         20'h0c181: data =  16'h0000; //               
         20'h0c182: data =  16'h0000; //               
         20'h0c183: data =  16'h0000; //               
         20'h0c184: data =  16'h7F80; //  11111111     
         20'h0c185: data =  16'h1DC0; //    111 111    
         20'h0c186: data =  16'h1CE0; //    111  111   
         20'h0c187: data =  16'h1CE0; //    111  111   
         20'h0c188: data =  16'h1CE0; //    111  111   
         20'h0c189: data =  16'h18E0; //    11   111   
         20'h0c18a: data =  16'h18E0; //    11   111   
         20'h0c18b: data =  16'h18C0; //    11   11    
         20'h0c18c: data =  16'h1980; //    11  11     
         20'h0c18d: data =  16'h1F00; //    11111      
         20'h0c18e: data =  16'h19C0; //    11  111    
         20'h0c18f: data =  16'h18C0; //    11   11    
         20'h0c190: data =  16'h18E0; //    11   111   
         20'h0c191: data =  16'h18E0; //    11   111   
         20'h0c192: data =  16'h18E0; //    11   111   
         20'h0c193: data =  16'h18E0; //    11   111   
         20'h0c194: data =  16'h30E0; //   11    111   
         20'h0c195: data =  16'h30E0; //   11    111   
         20'h0c196: data =  16'h31C0; //   11   111    
         20'h0c197: data =  16'h31C0; //   11   111    
         20'h0c198: data =  16'h3380; //   11  111     
         20'h0c199: data =  16'h7E00; //  111111       
         20'h0c19a: data =  16'h0000; //               
         20'h0c19b: data =  16'h0000; //               
         20'h0c19c: data =  16'h0000; //               
         20'h0c19d: data =  16'h0000; //               
         20'h0c19e: data =  16'h0000; //               
         20'h0c19f: data =  16'h0000; //
         
         /*C*/
         //code x0d1
         20'h0d1a0: data = 16'h0000; //               
         20'h0d1a1: data = 16'h0000; //               
         20'h0d1a2: data = 16'h0000; //               
         20'h0d1a3: data = 16'h0000; //               
         20'h0d1a4: data = 16'h0700; //      111      
         20'h0d1a5: data = 16'h0DE0; //     11 1111   
         20'h0d1a6: data = 16'h1DE0; //    111 1111   
         20'h0d1a7: data = 16'h1CE0; //    111  111   
         20'h0d1a8: data = 16'h1860; //    11    11   
         20'h0d1a9: data = 16'h1860; //    11    11   
         20'h0d1aa: data = 16'h3860; //   111    11   
         20'h0d1ab: data = 16'h3800; //   111         
         20'h0d1ac: data = 16'h3800; //   111         
         20'h0d1ad: data = 16'h3800; //   111         
         20'h0d1ae: data = 16'h3800; //   111         
         20'h0d1af: data = 16'h3800; //   111         
         20'h0d1b0: data = 16'h3800; //   111         
         20'h0d1b1: data = 16'h38E0; //   111   111   
         20'h0d1b2: data = 16'h38E0; //   111   111   
         20'h0d1b3: data = 16'h38E0; //   111   111   
         20'h0d1b4: data = 16'h38E0; //   111   111   
         20'h0d1b5: data = 16'h18C0; //    11   11    
         20'h0d1b6: data = 16'h18C0; //    11   11    
         20'h0d1b7: data = 16'h1DC0; //    111 111    
         20'h0d1b8: data = 16'h0D80; //     11 11     
         20'h0d1b9: data = 16'h0700; //      111      
         20'h0d1ba: data = 16'h0000; //               
         20'h0d1bb: data = 16'h0000; //               
         20'h0d1bc: data = 16'h0000; //               
         20'h0d1bd: data = 16'h0000; //               
         20'h0d1be: data = 16'h0000; //               
         20'h0d1bf: data = 16'h0000; //  
         
         /*D*/  
         //code x0e1
         20'h0e1c0: data = 16'h0000; //               
         20'h0e1c1: data = 16'h0000; //               
         20'h0e1c2: data = 16'h0000; //               
         20'h0e1c3: data = 16'h0000; //               
         20'h0e1c4: data = 16'h7F00; //  1111111      
         20'h0e1c5: data = 16'h1D80; //    111 11     
         20'h0e1c6: data = 16'h1DC0; //    111 111    
         20'h0e1c7: data = 16'h1CC0; //    111  11    
         20'h0e1c8: data = 16'h1CC0; //    111  11    
         20'h0e1c9: data = 16'h1CE0; //    111  111   
         20'h0e1ca: data = 16'h18E0; //    11   111   
         20'h0e1cb: data = 16'h18E0; //    11   111   
         20'h0e1cc: data = 16'h18E0; //    11   111   
         20'h0e1cd: data = 16'h18E0; //    11   111   
         20'h0e1ce: data = 16'h18E0; //    11   111   
         20'h0e1cf: data = 16'h18E0; //    11   111   
         20'h0e1d0: data = 16'h18E0; //    11   111   
         20'h0e1d1: data = 16'h18E0; //    11   111   
         20'h0e1d2: data = 16'h18C0; //    11   11    
         20'h0e1d3: data = 16'h19C0; //    11  111    
         20'h0e1d4: data = 16'h31C0; //   11   111    
         20'h0e1d5: data = 16'h3180; //   11   11     
         20'h0e1d6: data = 16'h3180; //   11   11     
         20'h0e1d7: data = 16'h3300; //   11  11      
         20'h0e1d8: data = 16'h3600; //   11 11       
         20'h0e1d9: data = 16'h7C00; //  11111        
         20'h0e1da: data = 16'h0000; //               
         20'h0e1db: data = 16'h0000; //               
         20'h0e1dc: data = 16'h0000; //               
         20'h0e1dd: data = 16'h0000; //               
         20'h0e1de: data = 16'h0000; //               
         20'h0e1df: data = 16'h0000; //               
         
         /*E*/
         //code x0f1
         20'h0f1e0: data = 16'h0000; //               
         20'h0f1e1: data = 16'h0000; //               
         20'h0f1e2: data = 16'h0000; //               
         20'h0f1e3: data = 16'h0000; //               
         20'h0f1e4: data = 16'h7FE0; //  1111111111   
         20'h0f1e5: data = 16'h1CC0; //    111  11    
         20'h0f1e6: data = 16'h1CC0; //    111  11    
         20'h0f1e7: data = 16'h1CC0; //    111  11    
         20'h0f1e8: data = 16'h1C00; //    111        
         20'h0f1e9: data = 16'h1C00; //    111        
         20'h0f1ea: data = 16'h1800; //    11         
         20'h0f1eb: data = 16'h1980; //    11  11     
         20'h0f1ec: data = 16'h1980; //    11  11     
         20'h0f1ed: data = 16'h1980; //    11  11     
         20'h0f1ee: data = 16'h1F80; //    111111     
         20'h0f1ef: data = 16'h1980; //    11  11     
         20'h0f1f0: data = 16'h1980; //    11  11     
         20'h0f1f1: data = 16'h1980; //    11  11     
         20'h0f1f2: data = 16'h1800; //    11         
         20'h0f1f3: data = 16'h1800; //    11         
         20'h0f1f4: data = 16'h3060; //   11     11   
         20'h0f1f5: data = 16'h3060; //   11     11   
         20'h0f1f6: data = 16'h3060; //   11     11   
         20'h0f1f7: data = 16'h3060; //   11     11   
         20'h0f1f8: data = 16'h3060; //   11     11   
         20'h0f1f9: data = 16'h7FE0; //  1111111111   
         20'h0f1fa: data = 16'h0000; //               
         20'h0f1fb: data = 16'h0000; //               
         20'h0f1fc: data = 16'h0000; //               
         20'h0f1fd: data = 16'h0000; //               
         20'h0f1fe: data = 16'h0000; //               
         20'h0f1ff: data = 16'h0000; //       
         
         /*F*/        
         //code x102
         20'h10200: data =16'h0000; //               
         20'h10201: data = 16'h0000; //               
         20'h10202: data = 16'h0000; //               
         20'h10203: data = 16'h0000; //               
         20'h10204: data = 16'h3FF8; //   11111111111 
         20'h10205: data = 16'h0E30; //     111   11  
         20'h10206: data = 16'h0E30; //     111   11  
         20'h10207: data = 16'h0E60; //     111  11   
         20'h10208: data = 16'h0E60; //     111  11   
         20'h10209: data = 16'h0E00; //     111       
         20'h1020a: data = 16'h0E00; //     111       
         20'h1020b: data = 16'h0EC0; //     111 11    
         20'h1020c: data = 16'h0EC0; //     111 11    
         20'h1020d: data = 16'h0EC0; //     111 11    
         20'h1020e: data = 16'h0FC0; //     111111    
         20'h1020f: data = 16'h0CC0; //     11  11    
         20'h10210: data = 16'h0CC0; //     11  11    
         20'h10211: data = 16'h0CC0; //     11  11    
         20'h10212: data = 16'h0C00; //     11        
         20'h10213: data = 16'h0C00; //     11        
         20'h10214: data = 16'h0C00; //     11        
         20'h10215: data = 16'h0C00; //     11        
         20'h10216: data = 16'h0C00; //     11        
         20'h10217: data = 16'h0C00; //     11        
         20'h10218: data = 16'h0C00; //     11        
         20'h10219: data = 16'h3C00; //   1111        
         20'h1021a: data = 16'h0000; //               
         20'h1021b: data = 16'h0000; //               
         20'h1021c: data = 16'h0000; //               
         20'h1021d: data = 16'h0000; //               
         20'h1021e: data = 16'h0000; //               
         20'h1021f: data = 16'h0000; //  
         
         /*G*/   
         //code x112
         20'h11220: data = 16'h0000; //               
         20'h11221: data = 16'h0000; //               
         20'h11222: data = 16'h0000; //               
         20'h11223: data = 16'h0000; //               
         20'h11224: data = 16'h0700; //      111      
         20'h11225: data = 16'h0DE0; //     11 1111   
         20'h11226: data = 16'h1DE0; //    111 1111   
         20'h11227: data = 16'h1CE0; //    111  111   
         20'h11228: data = 16'h1860; //    11    11   
         20'h11229: data = 16'h3860; //   111    11   
         20'h1122a: data = 16'h3860; //   111    11   
         20'h1122b: data = 16'h3860; //   111    11   
         20'h1122c: data = 16'h3800; //   111         
         20'h1122d: data = 16'h3800; //   111         
         20'h1122e: data = 16'h3800; //   111         
         20'h1122f: data = 16'h3BE0; //   111 11111   
         20'h11230: data = 16'h3BE0; //   111 11111   
         20'h11231: data = 16'h3EE0; //   11111 111   
         20'h11232: data = 16'h38E0; //   111   111   
         20'h11233: data = 16'h38E0; //   111   111   
         20'h11234: data = 16'h38E0; //   111   111   
         20'h11235: data = 16'h18C0; //    11   11    
         20'h11236: data = 16'h18C0; //    11   11    
         20'h11237: data = 16'h1DC0; //    111 111    
         20'h11238: data = 16'h0D80; //     11 11     
         20'h11239: data = 16'h0700; //      111      
         20'h1123a: data = 16'h0000; //               
         20'h1123b: data = 16'h0000; //               
         20'h1123c: data = 16'h0000; //               
         20'h1123d: data = 16'h0000; //               
         20'h1123e: data = 16'h0000; //               
         20'h1123f: data = 16'h0000; //  
         
         /*H*/
         //code x122
         20'h12240: data = 16'h0000; //               
         20'h12241: data = 16'h0000; //               
         20'h12242: data = 16'h0000; //               
         20'h12243: data = 16'h0000; //               
         20'h12244: data = 16'h7C78; //  11111   1111 
         20'h12245: data = 16'h1C60; //    111   11   
         20'h12246: data = 16'h1C60; //    111   11   
         20'h12247: data = 16'h1C60; //    111   11   
         20'h12248: data = 16'h1C60; //    111   11   
         20'h12249: data = 16'h1C60; //    111   11   
         20'h1224a: data = 16'h1C60; //    111   11   
         20'h1224b: data = 16'h1C60; //    111   11   
         20'h1224c: data = 16'h1C60; //    111   11   
         20'h1224d: data = 16'h1C60; //    111   11   
         20'h1224e: data = 16'h1FE0; //    11111111   
         20'h1224f: data = 16'h18E0; //    11   111   
         20'h12250: data = 16'h18E0; //    11   111   
         20'h12251: data = 16'h18E0; //    11   111   
         20'h12252: data = 16'h18E0; //    11   111   
         20'h12253: data = 16'h18E0; //    11   111   
         20'h12254: data = 16'h18E0; //    11   111   
         20'h12255: data = 16'h18E0; //    11   111   
         20'h12256: data = 16'h18E0; //    11   111   
         20'h12257: data = 16'h18E0; //    11   111   
         20'h12258: data = 16'h18E0; //    11   111   
         20'h12259: data = 16'h78F8; //  1111   11111 
         20'h1225a: data = 16'h0000; //               
         20'h1225b: data = 16'h0000; //               
         20'h1225c: data = 16'h0000; //               
         20'h1225d: data = 16'h0000; //               
         20'h1225e: data = 16'h0000; //               
         20'h1225f: data = 16'h0000; //  
         
         /*I*/
         //code x132
         20'h13260: data = 16'h0000; //               
         20'h13261: data = 16'h0000; //               
         20'h13262: data = 16'h0000; //               
         20'h13263: data = 16'h0000; //               
         20'h13264: data = 16'h1F80; //         
         20'h13265: data = 16'h0700; //          
         20'h13266: data = 16'h0700; //               
         20'h13267: data = 16'h0700; //    1111111    
         20'h13268: data = 16'h0700; //      111      
         20'h13269: data = 16'h0700; //      111      
         20'h1326a: data = 16'h0700; //      111      
         20'h1326b: data = 16'h0700; //      111      
         20'h1326c: data = 16'h0700; //      111      
         20'h1326d: data = 16'h0600; //      111      
         20'h1326e: data = 16'h0600; //      111      
         20'h1326f: data = 16'h0600; //      111      
         20'h13270: data = 16'h0600; //      111      
         20'h13271: data = 16'h0600; //      11       
         20'h13272: data = 16'h0600; //      11       
         20'h13273: data = 16'h0600; //      11       
         20'h13274: data = 16'h0600; //      11       
         20'h13275: data = 16'h0600; //      11       
         20'h13276: data = 16'h0600; //      11       
         20'h13277: data = 16'h0600; //      11       
         20'h13278: data = 16'h0600; //      11       
         20'h13279: data = 16'h1F80; //    111111     
         20'h1327a: data = 16'h0000; //               
         20'h1327b: data = 16'h0000; //               
         20'h1327c: data = 16'h0000; //               
         20'h1327d: data = 16'h0000; //               
         20'h1327e: data = 16'h0000; //               
         20'h1327f: data = 16'h0000; // 
         /*
         20'h13260: data = 16'h0000; //               
         20'h13261: data = 16'h0000; //               
         20'h13262: data = 16'h0000; //               
         20'h13263: data = 16'h0000; //               
         20'h13264: data = 16'h0F80; //     11111     
         20'h13265: data = 16'h0F80; //     11111     
         20'h13266: data = 16'h0000; //               
         20'h13267: data = 16'h1FC0; //    1111111    
         20'h13268: data = 16'h0700; //      111      
         20'h13269: data = 16'h0700; //      111      
         20'h1326a: data = 16'h0700; //      111      
         20'h1326b: data = 16'h0700; //      111      
         20'h1326c: data = 16'h0700; //      111      
         20'h1326d: data = 16'h0700; //      111      
         20'h1326e: data = 16'h0700; //      111      
         20'h1326f: data = 16'h0700; //      111      
         20'h13270: data = 16'h0700; //      111      
         20'h13271: data = 16'h0600; //      11       
         20'h13272: data = 16'h0600; //      11       
         20'h13273: data = 16'h0600; //      11       
         20'h13274: data = 16'h0600; //      11       
         20'h13275: data = 16'h0600; //      11       
         20'h13276: data = 16'h0600; //      11       
         20'h13277: data = 16'h0600; //      11       
         20'h13278: data = 16'h0600; //      11       
         20'h13279: data = 16'h1F80; //    111111     
         20'h1327a: data = 16'h0000; //               
         20'h1327b: data = 16'h0000; //               
         20'h1327c: data = 16'h0000; //               
         20'h1327d: data = 16'h0000; //               
         20'h1327e: data = 16'h0000; //               
         20'h1327f: data = 16'h0000; //  
         */ 
         
         /*J*/
         //code x142
         20'h14280: data = 16'h0000; //               
         20'h14281: data = 16'h0000; //               
         20'h14282: data = 16'h0000; //               
         20'h14283: data = 16'h0000; //               
         20'h14284: data = 16'h1FC0; //    1111111    
         20'h14285: data = 16'h0300; //       11      
         20'h14286: data = 16'h0300; //       11      
         20'h14287: data = 16'h0180; //        11     
         20'h14288: data = 16'h00C0; //         11    
         20'h14289: data = 16'h00C0; //         11    
         20'h1428a: data = 16'h00E0; //         111   
         20'h1428b: data = 16'h0060; //          11   
         20'h1428c: data = 16'h0070; //          111  
         20'h1428d: data = 16'h0070; //          111  
         20'h1428e: data = 16'h0070; //          111  
         20'h1428f: data = 16'h0070; //          111  
         20'h14290: data = 16'h3F70; //   111111 111  
         20'h14291: data = 16'h1870; //    11    111  
         20'h14292: data = 16'h3070; //   11     111  
         20'h14293: data = 16'h3070; //   11     111  
         20'h14294: data = 16'h3070; //   11     111  
         20'h14295: data = 16'h3060; //   11     11   
         20'h14296: data = 16'h30E0; //   11    111   
         20'h14297: data = 16'h38E0; //   111   111   
         20'h14298: data = 16'h19C0; //    11  111    
         20'h14299: data = 16'h0F80; //     11111     
         20'h1429a: data = 16'h0000; //               
         20'h1429b: data = 16'h0000; //               
         20'h1429c: data = 16'h0000; //               
         20'h1429d: data = 16'h0000; //               
         20'h1429e: data = 16'h0000; //               
         20'h1429f: data = 16'h0000; //      
         
         /*K*/
         //code x152
         20'h152a0: data = 16'h0000; //               
         20'h152a1: data = 16'h0000; //               
         20'h152a2: data = 16'h0000; //               
         20'h152a3: data = 16'h0000; //               
         20'h152a4: data = 16'h7DF0; //  11111 11111  
         20'h152a5: data = 16'h1CC0; //    111  11    
         20'h152a6: data = 16'h1CC0; //    111  11    
         20'h152a7: data = 16'h1D80; //    111 11     
         20'h152a8: data = 16'h1D80; //    111 11     
         20'h152a9: data = 16'h1F00; //    11111      
         20'h152aa: data = 16'h1F00; //    11111      
         20'h152ab: data = 16'h1E00; //    1111       
         20'h152ac: data = 16'h1E00; //    1111       
         20'h152ad: data = 16'h1E00; //    1111       
         20'h152ae: data = 16'h1E00; //    1111       
         20'h152af: data = 16'h1F00; //    11111      
         20'h152b0: data = 16'h1F00; //    11111      
         20'h152b1: data = 16'h1B00; //    11 11      
         20'h152b2: data = 16'h1B00; //    11 11      
         20'h152b3: data = 16'h1980; //    11  11     
         20'h152b4: data = 16'h1980; //    11  11     
         20'h152b5: data = 16'h1980; //    11  11     
         20'h152b6: data = 16'h18C0; //    11   11    
         20'h152b7: data = 16'h18C0; //    11   11    
         20'h152b8: data = 16'h18C0; //    11   11    
         20'h152b9: data = 16'h79F0; //  1111  11111  
         20'h152ba: data = 16'h0000; //               
         20'h152bb: data = 16'h0000; //               
         20'h152bc: data = 16'h0000; //               
         20'h152bd: data = 16'h0000; //               
         20'h152be: data = 16'h0000; //               
         20'h152bf: data = 16'h0000; //              
         
         /*L*/ 
         //code x162
         20'h162c0: data = 16'h0000; //               
         20'h162c1: data = 16'h0000; //               
         20'h162c2: data = 16'h0000; //               
         20'h162c3: data = 16'h0000; //               
         20'h162c4: data = 16'h3E00; //   11111       
         20'h162c5: data = 16'h0E00; //     111       
         20'h162c6: data = 16'h0E00; //     111       
         20'h162c7: data = 16'h0E00; //     111       
         20'h162c8: data = 16'h0E00; //     111       
         20'h162c9: data = 16'h0E00; //     111       
         20'h162ca: data = 16'h0E00; //     111       
         20'h162cb: data = 16'h0E00; //     111       
         20'h162cc: data = 16'h0E00; //     111       
         20'h162cd: data = 16'h0E00; //     111       
         20'h162ce: data = 16'h0E00; //     111       
         20'h162cf: data = 16'h0C00; //     11        
         20'h162d0: data = 16'h0C00; //     11        
         20'h162d1: data = 16'h0C00; //     11        
         20'h162d2: data = 16'h0C60; //     11   11   
         20'h162d3: data = 16'h0C60; //     11   11   
         20'h162d4: data = 16'h0C60; //     11   11   
         20'h162d5: data = 16'h0C60; //     11   11   
         20'h162d6: data = 16'h0C60; //     11   11   
         20'h162d7: data = 16'h0C60; //     11   11   
         20'h162d8: data = 16'h0C60; //     11   11   
         20'h162d9: data = 16'h3FE0; //   111111111   
         20'h162da: data = 16'h0000; //               
         20'h162db: data = 16'h0000; //               
         20'h162dc: data = 16'h0000; //               
         20'h162dd: data = 16'h0000; //               
         20'h162de: data = 16'h0000; //               
         20'h162df: data = 16'h0000; //   
               
         /*M*/    
         //code x172
         20'h172e0: data = 16'h0000; //               
         20'h172e1: data = 16'h0000; //               
         20'h172e2: data = 16'h0000; //               
         20'h172e3: data = 16'h0000; //               
         20'h172e4: data = 16'hF83C; // 11111     1111
         20'h172e5: data = 16'h3C30; //   1111    11  
         20'h172e6: data = 16'h3C70; //   1111   111  
         20'h172e7: data = 16'h3C70; //   1111   111  
         20'h172e8: data = 16'h3C70; //   1111   111  
         20'h172e9: data = 16'h3CF0; //   1111  1111  
         20'h172ea: data = 16'h3EF0; //   11111 1111  
         20'h172eb: data = 16'h3EF0; //   11111 1111  
         20'h172ec: data = 16'h3FB0; //   1111111 11  
         20'h172ed: data = 16'h3FB0; //   1111111 11  
         20'h172ee: data = 16'h3BB0; //   111 111 11  
         20'h172ef: data = 16'h3BB0; //   111 111 11  
         20'h172f0: data = 16'h3330; //   11  11  11  
         20'h172f1: data = 16'h3370; //   11  11 111  
         20'h172f2: data = 16'h3370; //   11  11 111  
         20'h172f3: data = 16'h3070; //   11     111  
         20'h172f4: data = 16'h3070; //   11     111  
         20'h172f5: data = 16'h3070; //   11     111  
         20'h172f6: data = 16'h3070; //   11     111  
         20'h172f7: data = 16'h3070; //   11     111  
         20'h172f8: data = 16'h3070; //   11     111  
         20'h172f9: data = 16'hF07C; // 1111     11111
         20'h172fa: data = 16'h0000; //               
         20'h172fb: data = 16'h0000; //               
         20'h172fc: data = 16'h0000; //               
         20'h172fd: data = 16'h0000; //               
         20'h172fe: data = 16'h0000; //               
         20'h172ff: data = 16'h0000; // 
         
         /*N*/             
         //code x183
         20'h18300: data = 16'h0000; //               
         20'h18301: data = 16'h0000; //               
         20'h18302: data = 16'h0000; //               
         20'h18303: data = 16'h0000; //               
         20'h18304: data = 16'h7C78; //  11111   1111 
         20'h18305: data = 16'h1C60; //    111   11   
         20'h18306: data = 16'h1E60; //    1111  11   
         20'h18307: data = 16'h1E60; //    1111  11   
         20'h18308: data = 16'h1E60; //    1111  11   
         20'h18309: data = 16'h1E60; //    1111  11   
         20'h1830a: data = 16'h1E60; //    1111  11   
         20'h1830b: data = 16'h1E60; //    1111  11   
         20'h1830c: data = 16'h1E60; //    1111  11   
         20'h1830d: data = 16'h1F60; //    11111 11   
         20'h1830e: data = 16'h1FE0; //    11111111   
         20'h1830f: data = 16'h1FE0; //    11111111   
         20'h18310: data = 16'h1BE0; //    11 11111   
         20'h18311: data = 16'h1BE0; //    11 11111   
         20'h18312: data = 16'h1BE0; //    11 11111   
         20'h18313: data = 16'h1BE0; //    11 11111   
         20'h18314: data = 16'h19E0; //    11  1111   
         20'h18315: data = 16'h19E0; //    11  1111   
         20'h18316: data = 16'h19E0; //    11  1111   
         20'h18317: data = 16'h19E0; //    11  1111   
         20'h18318: data = 16'h18E0; //    11   111   
         20'h18319: data = 16'h78F8; //  1111   11111 
         20'h1831a: data = 16'h0000; //               
         20'h1831b: data = 16'h0000; //               
         20'h1831c: data = 16'h0000; //               
         20'h1831d: data = 16'h0000; //               
         20'h1831e: data = 16'h0000; //               
         20'h1831f: data = 16'h0000; //  
         
         /*O*/
         //code x193
         20'h19320: data = 16'h0000; //               
         20'h19321: data = 16'h0000; //               
         20'h19322: data = 16'h0000; //               
         20'h19323: data = 16'h0000; //               
         20'h19324: data = 16'h0780; //      1111     
         20'h19325: data = 16'h0CC0; //     11  11    
         20'h19326: data = 16'h1CE0; //    111  111   
         20'h19327: data = 16'h1860; //    11    11   
         20'h19328: data = 16'h1860; //    11    11   
         20'h19329: data = 16'h3870; //   111    111  
         20'h1932a: data = 16'h3870; //   111    111  
         20'h1932b: data = 16'h3870; //   111    111  
         20'h1932c: data = 16'h3870; //   111    111  
         20'h1932d: data = 16'h3870; //   111    111  
         20'h1932e: data = 16'h3870; //   111    111  
         20'h1932f: data = 16'h3870; //   111    111  
         20'h19330: data = 16'h3870; //   111    111  
         20'h19331: data = 16'h3870; //   111    111  
         20'h19332: data = 16'h3870; //   111    111  
         20'h19333: data = 16'h3870; //   111    111  
         20'h19334: data = 16'h3870; //   111    111  
         20'h19335: data = 16'h1860; //    11    11   
         20'h19336: data = 16'h1860; //    11    11   
         20'h19337: data = 16'h1CE0; //    111  111   
         20'h19338: data = 16'h0CC0; //     11  11    
         20'h19339: data = 16'h0780; //      1111     
         20'h1933a: data = 16'h0000; //               
         20'h1933b: data = 16'h0000; //               
         20'h1933c: data = 16'h0000; //               
         20'h1933d: data = 16'h0000; //               
         20'h1933e: data = 16'h0000; //               
         20'h1933f: data = 16'h0000; // 
         
         /*P*/
         //code x1a3
         20'h1a340: data = 16'h0000; //               
         20'h1a341: data = 16'h0000; //               
         20'h1a342: data = 16'h0000; //               
         20'h1a343: data = 16'h0000; //               
         20'h1a344: data = 16'h3F80; //   1111111     
         20'h1a345: data = 16'h0EC0; //     111 11    
         20'h1a346: data = 16'h0EE0; //     111 111   
         20'h1a347: data = 16'h0E70; //     111  111  
         20'h1a348: data = 16'h0E70; //     111  111  
         20'h1a349: data = 16'h0E70; //     111  111  
         20'h1a34a: data = 16'h0E70; //     111  111  
         20'h1a34b: data = 16'h0E70; //     111  111  
         20'h1a34c: data = 16'h0E70; //     111  111  
         20'h1a34d: data = 16'h0EE0; //     111 111   
         20'h1a34e: data = 16'h0EE0; //     111 111   
         20'h1a34f: data = 16'h0DC0; //     11 111    
         20'h1a350: data = 16'h0F80; //     11111     
         20'h1a351: data = 16'h0C00; //     11        
         20'h1a352: data = 16'h0C00; //     11        
         20'h1a353: data = 16'h0C00; //     11        
         20'h1a354: data = 16'h0C00; //     11        
         20'h1a355: data = 16'h0C00; //     11        
         20'h1a356: data = 16'h0C00; //     11        
         20'h1a357: data = 16'h0C00; //     11        
         20'h1a358: data = 16'h0C00; //     11        
         20'h1a359: data = 16'h3C00; //   1111        
         20'h1a35a: data = 16'h0000; //               
         20'h1a35b: data = 16'h0000; //               
         20'h1a35c: data = 16'h0000; //               
         20'h1a35d: data = 16'h0000; //               
         20'h1a35e: data = 16'h0000; //               
         20'h1a35f: data = 16'h0000; //  
         
         /*Q*/       
         //code x1b3
         20'h1b360: data = 16'h0000; //               
         20'h1b361: data = 16'h0000; //               
         20'h1b362: data = 16'h0000; //               
         20'h1b363: data = 16'h0000; //               
         20'h1b364: data = 16'h0780; //      1111     
         20'h1b365: data = 16'h0CC0; //     11  11    
         20'h1b366: data = 16'h1CE0; //    111  111   
         20'h1b367: data = 16'h1860; //    11    11   
         20'h1b368: data = 16'h1860; //    11    11   
         20'h1b369: data = 16'h3870; //   111    111  
         20'h1b36a: data = 16'h3870; //   111    111  
         20'h1b36b: data = 16'h3870; //   111    111  
         20'h1b36c: data = 16'h3870; //   111    111  
         20'h1b36d: data = 16'h3870; //   111    111  
         20'h1b36e: data = 16'h3870; //   111    111  
         20'h1b36f: data = 16'h3870; //   111    111  
         20'h1b370: data = 16'h3870; //   111    111  
         20'h1b371: data = 16'h3870; //   111    111  
         20'h1b372: data = 16'h3870; //   111    111  
         20'h1b373: data = 16'h3870; //   111    111  
         20'h1b374: data = 16'h3860; //   111    11   
         20'h1b375: data = 16'h1FE0; //    11111111   
         20'h1b376: data = 16'h1B60; //    11 11 11   
         20'h1b377: data = 16'h1FC0; //    1111111    
         20'h1b378: data = 16'h0DC0; //     11 111    
         20'h1b379: data = 16'h0780; //      1111     
         20'h1b37a: data = 16'h00C0; //         11    
         20'h1b37b: data = 16'h00C0; //         11    
         20'h1b37c: data = 16'h0060; //          11   
         20'h1b37d: data = 16'h01F0; //        11111  
         20'h1b37e: data = 16'h0000; //               
         20'h1b37f: data = 16'h0000; //     
                
         /*R*/
         //code x1c3
         20'h1c380: data = 16'h0000; //               
         20'h1c381: data = 16'h0000; //               
         20'h1c382: data = 16'h0000; //               
         20'h1c383: data = 16'h0000; //               
         20'h1c384: data = 16'h7F00; //  1111111      
         20'h1c385: data = 16'h1D80; //    111 11     
         20'h1c386: data = 16'h1DC0; //    111 111    
         20'h1c387: data = 16'h1CE0; //    111  111   
         20'h1c388: data = 16'h1CE0; //    111  111   
         20'h1c389: data = 16'h1CE0; //    111  111   
         20'h1c38a: data = 16'h1CE0; //    111  111   
         20'h1c38b: data = 16'h1CE0; //    111  111   
         20'h1c38c: data = 16'h1CE0; //    111  111   
         20'h1c38d: data = 16'h1DC0; //    111 111    
         20'h1c38e: data = 16'h1DC0; //    111 111    
         20'h1c38f: data = 16'h1B80; //    11 111     
         20'h1c390: data = 16'h1E00; //    1111       
         20'h1c391: data = 16'h1E00; //    1111       
         20'h1c392: data = 16'h1F00; //    11111      
         20'h1c393: data = 16'h1B00; //    11 11      
         20'h1c394: data = 16'h1B00; //    11 11      
         20'h1c395: data = 16'h1980; //    11  11     
         20'h1c396: data = 16'h1980; //    11  11     
         20'h1c397: data = 16'h18C0; //    11   11    
         20'h1c398: data = 16'h18C0; //    11   11    
         20'h1c399: data = 16'h7BF0; //  1111 111111  
         20'h1c39a: data = 16'h0000; //               
         20'h1c39b: data = 16'h0000; //               
         20'h1c39c: data = 16'h0000; //               
         20'h1c39d: data = 16'h0000; //               
         20'h1c39e: data = 16'h0000; //               
         20'h1c39f: data = 16'h0000; //    
         
         /*S*/  
         //code x1d3
         20'h1d3a0: data = 16'h0000; //               
         20'h1d3a1: data = 16'h0000; //               
         20'h1d3a2: data = 16'h0000; //               
         20'h1d3a3: data = 16'h0000; //               
         20'h1d3a4: data = 16'h0FC0; //     111111    
         20'h1d3a5: data = 16'h1FC0; //    1111111    
         20'h1d3a6: data = 16'h39C0; //   111  111    
         20'h1d3a7: data = 16'h38C0; //   111   11    
         20'h1d3a8: data = 16'h38C0; //   111   11    
         20'h1d3a9: data = 16'h38C0; //   111   11    
         20'h1d3aa: data = 16'h38C0; //   111   11    
         20'h1d3ab: data = 16'h1800; //    11         
         20'h1d3ac: data = 16'h1C00; //    111        
         20'h1d3ad: data = 16'h0E00; //     111       
         20'h1d3ae: data = 16'h0600; //      11       
         20'h1d3af: data = 16'h0300; //       11      
         20'h1d3b0: data = 16'h0180; //        11     
         20'h1d3b1: data = 16'h61C0; //  11    111    
         20'h1d3b2: data = 16'h61C0; //  11    111    
         20'h1d3b3: data = 16'h61C0; //  11    111    
         20'h1d3b4: data = 16'h61C0; //  11    111    
         20'h1d3b5: data = 16'h61C0; //  11    111    
         20'h1d3b6: data = 16'h71C0; //  111   111    
         20'h1d3b7: data = 16'h7180; //  111   11     
         20'h1d3b8: data = 16'h7B80; //  1111 111     
         20'h1d3b9: data = 16'h0F00; //     1111      
         20'h1d3ba: data = 16'h0000; //               
         20'h1d3bb: data = 16'h0000; //               
         20'h1d3bc: data = 16'h0000; //               
         20'h1d3bd: data = 16'h0000; //               
         20'h1d3be: data = 16'h0000; //               
         20'h1d3bf: data = 16'h0000; //  
         
         /*T*/
         //code x1e3
         20'h1e3c0: data = 16'h0000; //               
         20'h1e3c1: data = 16'h0000; //               
         20'h1e3c2: data = 16'h0000; //               
         20'h1e3c3: data = 16'h0000; //               
         20'h1e3c4: data = 16'h3FF0; //   1111111111  
         20'h1e3c5: data = 16'h3370; //   11  11 111  
         20'h1e3c6: data = 16'h3330; //   11  11  11  
         20'h1e3c7: data = 16'h3330; //   11  11  11  
         20'h1e3c8: data = 16'h3330; //   11  11  11  
         20'h1e3c9: data = 16'h3330; //   11  11  11  
         20'h1e3ca: data = 16'h3330; //   11  11  11  
         20'h1e3cb: data = 16'h3330; //   11  11  11  
         20'h1e3cc: data = 16'h0300; //       11      
         20'h1e3cd: data = 16'h0300; //       11      
         20'h1e3ce: data = 16'h0300; //       11      
         20'h1e3cf: data = 16'h0700; //      111      
         20'h1e3d0: data = 16'h0700; //      111      
         20'h1e3d1: data = 16'h0700; //      111      
         20'h1e3d2: data = 16'h0700; //      111      
         20'h1e3d3: data = 16'h0700; //      111      
         20'h1e3d4: data = 16'h0700; //      111      
         20'h1e3d5: data = 16'h0700; //      111      
         20'h1e3d6: data = 16'h0700; //      111      
         20'h1e3d7: data = 16'h0700; //      111      
         20'h1e3d8: data = 16'h0700; //      111      
         20'h1e3d9: data = 16'h1FC0; //    1111111    
         20'h1e3da: data = 16'h0000; //               
         20'h1e3db: data = 16'h0000; //               
         20'h1e3dc: data = 16'h0000; //               
         20'h1e3dd: data = 16'h0000; //               
         20'h1e3de: data = 16'h0000; //               
         20'h1e3df: data = 16'h0000; //    
         
         /*U*/     
         //code x1f3        
         20'h1f3e0: data = 16'h0000; //               
         20'h1f3e1: data = 16'h0000; //               
         20'h1f3e2: data = 16'h0000; //               
         20'h1f3e3: data = 16'h0000; //               
         20'h1f3e4: data = 16'h1F00; //    11111      
         20'h1f3e5: data = 16'h0C00; //     11        
         20'h1f3e6: data = 16'h0FF0; //     11111111  
         20'h1f3e7: data = 16'h0CC0; //     11  11    
         20'h1f3e8: data = 16'h0CC0; //     11  11    
         20'h1f3e9: data = 16'h1860; //    11    11   
         20'h1f3ea: data = 16'h1860; //    11    11   
         20'h1f3eb: data = 16'h1870; //    11    111  
         20'h1f3ec: data = 16'h1870; //    11    111  
         20'h1f3ed: data = 16'h3870; //   111    111  
         20'h1f3ee: data = 16'h3870; //   111    111  
         20'h1f3ef: data = 16'h3870; //   111    111  
         20'h1f3f0: data = 16'h3870; //   111    111  
         20'h1f3f1: data = 16'h3870; //   111    111  
         20'h1f3f2: data = 16'h3870; //   111    111  
         20'h1f3f3: data = 16'h3860; //   111    11   
         20'h1f3f4: data = 16'h38E0; //   111   111   
         20'h1f3f5: data = 16'h38E0; //   111   111   
         20'h1f3f6: data = 16'h18C0; //    11   11    
         20'h1f3f7: data = 16'h1CC0; //    111  11    
         20'h1f3f8: data = 16'h0D80; //     11 11     
         20'h1f3f9: data = 16'h0700; //      111      
         20'h1f3fa: data = 16'h0000; //               
         20'h1f3fb: data = 16'h0000; //               
         20'h1f3fc: data = 16'h0000; //               
         20'h1f3fd: data = 16'h0000; //               
         20'h1f3fe: data = 16'h0000; //               
         20'h1f3ff: data = 16'h0000; //  
                    
         /*V*/
        //code x204
         20'h20400: data = 16'h0000; //               
         20'h20401: data = 16'h0000; //               
         20'h20402: data = 16'h0000; //               
         20'h20403: data = 16'h0000; //               
         20'h20404: data = 16'h7CF8; //  11111  11111 
         20'h20405: data = 16'h1C60; //    111   11   
         20'h20406: data = 16'h1C60; //    111   11   
         20'h20407: data = 16'h1C60; //    111   11   
         20'h20408: data = 16'h1C60; //    111   11   
         20'h20409: data = 16'h1CC0; //    111  11    
         20'h2040a: data = 16'h0CC0; //     11  11    
         20'h2040b: data = 16'h0CC0; //     11  11    
         20'h2040c: data = 16'h0CC0; //     11  11    
         20'h2040d: data = 16'h0EC0; //     111 11    
         20'h2040e: data = 16'h0EC0; //     111 11    
         20'h2040f: data = 16'h0F80; //     11111     
         20'h20410: data = 16'h0780; //      1111     
         20'h20411: data = 16'h0780; //      1111     
         20'h20412: data = 16'h0780; //      1111     
         20'h20413: data = 16'h0780; //      1111     
         20'h20414: data = 16'h0780; //      1111     
         20'h20415: data = 16'h0700; //      111      
         20'h20416: data = 16'h0700; //      111      
         20'h20417: data = 16'h0300; //       11      
         20'h20418: data = 16'h0300; //       11      
         20'h20419: data = 16'h0700; //      111      
         20'h2041a: data = 16'h0000; //               
         20'h2041b: data = 16'h0000; //               
         20'h2041c: data = 16'h0000; //               
         20'h2041d: data = 16'h0000; //               
         20'h2041e: data = 16'h0000; //               
         20'h2041f: data = 16'h0000; // 
            
         /*W*/ 
         //code x214
         20'h21420: data = 16'h0000; //               
         20'h21421: data = 16'h0000; //               
         20'h21422: data = 16'h0000; //               
         20'h21423: data = 16'h0000; //               
         20'h21424: data = 16'hF83C; // 11111     1111
         20'h21425: data = 16'h3830; //   111     11  
         20'h21426: data = 16'h3830; //   111     11  
         20'h21427: data = 16'h3830; //   111     11  
         20'h21428: data = 16'h3830; //   111     11  
         20'h21429: data = 16'h3830; //   111     11  
         20'h2142a: data = 16'h3830; //   111     11  
         20'h2142b: data = 16'h3B30; //   111 11  11  
         20'h2142c: data = 16'h3B30; //   111 11  11  
         20'h2142d: data = 16'h3330; //   11  11  11  
         20'h2142e: data = 16'h3770; //   11 111 111  
         20'h2142f: data = 16'h3770; //   11 111 111  
         20'h21430: data = 16'h37F0; //   11 1111111  
         20'h21431: data = 16'h37F0; //   11 1111111  
         20'h21432: data = 16'h3DF0; //   1111 11111  
         20'h21433: data = 16'h3DF0; //   1111 11111  
         20'h21434: data = 16'h3DF0; //   1111 11111  
         20'h21435: data = 16'h39F0; //   111  11111  
         20'h21436: data = 16'h38F0; //   111   1111  
         20'h21437: data = 16'h38F0; //   111   1111  
         20'h21438: data = 16'h30F0; //   11    1111  
         20'h21439: data = 16'hF07C; // 1111     11111
         20'h2143a: data = 16'h0000; //               
         20'h2143b: data = 16'h0000; //               
         20'h2143c: data = 16'h0000; //               
         20'h2143d: data = 16'h0000; //               
         20'h2143e: data = 16'h0000; //               
         20'h2143f: data = 16'h0000; //  
         
         /*X*/   
         //code x224
         20'h22440: data = 16'h0000; //               
         20'h22441: data = 16'h0000; //               
         20'h22442: data = 16'h0000; //               
         20'h22443: data = 16'h0000; //               
         20'h22444: data = 16'h7DF8; //  11111 111111 
         20'h22445: data = 16'h1860; //    11    11   
         20'h22446: data = 16'h18C0; //    11   11    
         20'h22447: data = 16'h18C0; //    11   11    
         20'h22448: data = 16'h0CC0; //     11  11    
         20'h22449: data = 16'h0D80; //     11 11     
         20'h2244a: data = 16'h0D80; //     11 11     
         20'h2244b: data = 16'h0780; //      1111     
         20'h2244c: data = 16'h0700; //      111      
         20'h2244d: data = 16'h0700; //      111      
         20'h2244e: data = 16'h0700; //      111      
         20'h2244f: data = 16'h0300; //       11      
         20'h22450: data = 16'h0700; //      111      
         20'h22451: data = 16'h0780; //      1111     
         20'h22452: data = 16'h0F80; //     11111     
         20'h22453: data = 16'h0D80; //     11 11     
         20'h22454: data = 16'h0DC0; //     11 111    
         20'h22455: data = 16'h19C0; //    11  111    
         20'h22456: data = 16'h18E0; //    11   111   
         20'h22457: data = 16'h18E0; //    11   111   
         20'h22458: data = 16'h30E0; //   11    111   
         20'h22459: data = 16'h7CF8; //  11111  11111 
         20'h2245a: data = 16'h0000; //               
         20'h2245b: data = 16'h0000; //               
         20'h2245c: data = 16'h0000; //               
         20'h2245d: data = 16'h0000; //               
         20'h2245e: data = 16'h0000; //               
         20'h2245f: data = 16'h0000; // 
          
         /*Y*/             
         //code x234
         20'h23460: data = 16'h0000; //               
         20'h23461: data = 16'h0000; //               
         20'h23462: data = 16'h0000; //               
         20'h23463: data = 16'h0000; //               
         20'h23464: data = 16'h7EF8; //  111111 11111 
         20'h23465: data = 16'h1860; //    11    11   
         20'h23466: data = 16'h1860; //    11    11   
         20'h23467: data = 16'h1C60; //    111   11   
         20'h23468: data = 16'h0C60; //     11   11   
         20'h23469: data = 16'h0EC0; //     111 11    
         20'h2346a: data = 16'h0EC0; //     111 11    
         20'h2346b: data = 16'h07C0; //      11111    
         20'h2346c: data = 16'h0780; //      1111     
         20'h2346d: data = 16'h0780; //      1111     
         20'h2346e: data = 16'h0780; //      1111     
         20'h2346f: data = 16'h0300; //       11      
         20'h23470: data = 16'h0300; //       11      
         20'h23471: data = 16'h0300; //       11      
         20'h23472: data = 16'h0300; //       11      
         20'h23473: data = 16'h0300; //       11      
         20'h23474: data = 16'h0300; //       11      
         20'h23475: data = 16'h0380; //       111     
         20'h23476: data = 16'h0380; //       111     
         20'h23477: data = 16'h0380; //       111     
         20'h23478: data = 16'h0380; //       111     
         20'h23479: data = 16'h0FC0; //     111111    
         20'h2347a: data = 16'h0000; //               
         20'h2347b: data = 16'h0000; //               
         20'h2347c: data = 16'h0000; //               
         20'h2347d: data = 16'h0000; //               
         20'h2347e: data = 16'h0000; //               
         20'h2347f: data = 16'h0000; // 
         
         /*Z*/
         //code x244
         20'h24480: data = 16'h0000; //               
         20'h24481: data = 16'h0000; //               
         20'h24482: data = 16'h0000; //               
         20'h24483: data = 16'h0000; //               
         20'h24484: data = 16'h1FF0; //    111111111  
         20'h24485: data = 16'h18E0; //    11   111   
         20'h24486: data = 16'h18E0; //    11   111   
         20'h24487: data = 16'h18E0; //    11   111   
         20'h24488: data = 16'h19C0; //    11  111    
         20'h24489: data = 16'h19C0; //    11  111    
         20'h2448a: data = 16'h31C0; //   11   111    
         20'h2448b: data = 16'h3180; //   11   11     
         20'h2448c: data = 16'h0380; //       111     
         20'h2448d: data = 16'h0300; //       11      
         20'h2448e: data = 16'h0300; //       11      
         20'h2448f: data = 16'h0700; //      111      
         20'h24490: data = 16'h0600; //      11       
         20'h24491: data = 16'h0600; //      11       
         20'h24492: data = 16'h0E60; //     111  11   
         20'h24493: data = 16'h0C60; //     11   11   
         20'h24494: data = 16'h0C60; //     11   11   
         20'h24495: data = 16'h1860; //    11    11   
         20'h24496: data = 16'h1860; //    11    11   
         20'h24497: data = 16'h1860; //    11    11   
         20'h24498: data = 16'h3060; //   11     11   
         20'h24499: data = 16'h3FE0; //   111111111   
         20'h2449a: data = 16'h0000; //               
         20'h2449b: data = 16'h0000; //               
         20'h2449c: data = 16'h0000; //               
         20'h2449d: data = 16'h0000; //               
         20'h2449e: data = 16'h0000; //               
         20'h2449f: data = 16'h0000; //
         
         default:   data = 16'h0000;
         /*               
         //code x25   
         20'h004a0: data = 8'b00000000; // 
         20'h004a1: data = 8'b00000000; // 
         20'h004a2: data = 8'b00011100; //    ****
         20'h004a3: data = 8'b00001100; //     **
         20'h004a4: data = 8'b00001100; //     **
         20'h004a5: data = 8'b00001100; //     **
         20'h004a6: data = 8'b00001100; //     **
         20'h004a7: data = 8'b00001100; //     **
         20'h004a8: data = 8'b01001100; // **  **
         20'h004a9: data = 8'b01001100; // **  **
         20'h004aa: data = 8'b01001100; // **  **
         20'h004ab: data = 8'b01111000; //  ****
         20'h004ac: data = 8'b00000000; // 
         20'h004ad: data = 8'b00000000; // 
         20'h004ae: data = 8'b00000000; // 
         20'h004af: data = 8'b00000000; //    
         20'h004b0: data = 8'b00000000; // 
         20'h004b1: data = 8'b00000000; // 
         20'h004b2: data = 8'b01100100; // ***  **
         20'h004b3: data = 8'b01100100; //  **  **
         20'h004b4: data = 8'b01100100; //  **  **
         20'h004b5: data = 8'b01101100; //  ** **
         20'h004b6: data = 8'b01111000; //  ****
         20'h004b7: data = 8'b01111000; //  ****
         20'h004b8: data = 8'b01101100; //  ** **
         20'h004b9: data = 8'b01100100; //  **  **
         20'h004ba: data = 8'b01100100; //  **  **
         20'h004bb: data = 8'b01100100; // ***  **
         20'h004bc: data = 8'b00000000; // 
         20'h004bd: data = 8'b00000000; // 
         20'h004be: data = 8'b00000000; // 
         20'h004bf: data = 8'b00000000; // 
         
         //code x4c   
         20'h004c0: data = 8'b00000000; // 
         20'h004c1: data = 8'b00000000; // 
         20'h004c2: data = 8'b01110000; // ****
         20'h004c3: data = 8'b01100000; //  **
         20'h004c4: data = 8'b01100000; //  **
         20'h004c5: data = 8'b01100000; //  **
         20'h004c6: data = 8'b01100000; //  **
         20'h004c7: data = 8'b01100000; //  **
         20'h004c8: data = 8'b01100000; //  **
         20'h004c9: data = 8'b01100000; //  **   *
         20'h004ca: data = 8'b01100100; //  **  **
         20'h004cb: data = 8'b01111100; // *******
         20'h004cc: data = 8'b00000000; // 
         20'h004cd: data = 8'b00000000; // 
         20'h004ce: data = 8'b00000000; // 
         20'h004cf: data = 8'b00000000; // 
         //code x4d   
         20'h004d0: data = 8'b00000000; // 
         20'h004d1: data = 8'b00000000; // 
         20'h004d2: data = 8'b01000010; // **    **
         20'h004d3: data = 8'b01100110; // ***  ***
         20'h004d4: data = 8'b01111110; // ********
         20'h004d5: data = 8'b01111110; // ********
         20'h004d6: data = 8'b01011010; // ** ** **
         20'h004d7: data = 8'b01000010; // **    **
         20'h004d8: data = 8'b01000010; // **    **
         20'h004d9: data = 8'b01000010; // **    **
         20'h004da: data = 8'b01000010; // **    **
         20'h004db: data = 8'b01000010; // **    **
         20'h004dc: data = 8'b00000000; // 
         20'h004dd: data = 8'b00000000; // 
         20'h004de: data = 8'b00000000; // 
         20'h004df: data = 8'b00000000; // 
         //code x4e   
         20'h004e0: data = 8'b00000000; // 
         20'h004e1: data = 8'b00000000; // 
         20'h004e2: data = 8'b01000100; // **   **
         20'h004e3: data = 8'b01100100; // ***  **
         20'h004e4: data = 8'b01110100; // **** **
         20'h004e5: data = 8'b01111100; // *******
         20'h004e6: data = 8'b01011100; // ** ****
         20'h004e7: data = 8'b01001100; // **  ***
         20'h004e8: data = 8'b01000100; // **   **
         20'h004e9: data = 8'b01000100; // **   **
         20'h004ea: data = 8'b01000100; // **   **
         20'h004eb: data = 8'b01000100; // **   **
         20'h004ec: data = 8'b00000000; // 
         20'h004ed: data = 8'b00000000; // 
         20'h004ee: data = 8'b00000000; // 
         20'h004ef: data = 8'b00000000; // 
         //code x4f   
         20'h004f0: data = 8'b00000000; // 
         20'h004f1: data = 8'b00000000; // 
         20'h004f2: data = 8'b01111100; //  *****
         20'h004f3: data = 8'b01000100; // **   **
         20'h004f4: data = 8'b01000100; // **   **
         20'h004f5: data = 8'b01000100; // **   **
         20'h004f6: data = 8'b01000100; // **   **
         20'h004f7: data = 8'b01000100; // **   **
         20'h004f8: data = 8'b01000100; // **   **
         20'h004f9: data = 8'b01000100; // **   **
         20'h004fa: data = 8'b01000100; // **   **
         20'h004fb: data = 8'b01111100; //  *****
         20'h004fc: data = 8'b00000000; // 
         20'h004fd: data = 8'b00000000; // 
         20'h004fe: data = 8'b00000000; // 
         20'h004ff: data = 8'b00000000; // 
         //code x50   
         20'h00500: data = 8'b00000000; // 
         20'h00501: data = 8'b00000000; // 
         20'h00502: data = 8'b01111100; // ******
         20'h00503: data = 8'b01100100; //  **  **
         20'h00504: data = 8'b01100100; //  **  **
         20'h00505: data = 8'b01100100; //  **  **
         20'h00506: data = 8'b01111100; //  *****
         20'h00507: data = 8'b01100000; //  **
         20'h00508: data = 8'b01100000; //  **
         20'h00509: data = 8'b01100000; //  **
         20'h0050a: data = 8'b01100000; //  **
         20'h0050b: data = 8'b01110000; // ****
         20'h0050c: data = 8'b00000000; // 
         20'h0050d: data = 8'b00000000; // 
         20'h0050e: data = 8'b00000000; // 
         20'h0050f: data = 8'b00000000; // 
         //code x51
         20'h00510: data = 8'b00000000; // 
         20'h00511: data = 8'b00000000; // 
         20'h00512: data = 8'b01111100; //  *****
         20'h00513: data = 8'b01000100; // **   **
         20'h00514: data = 8'b01000100; // **   **
         20'h00515: data = 8'b01000100; // **   **
         20'h00516: data = 8'b01000100; // **   **
         20'h00517: data = 8'b01000100; // **   **
         20'h00518: data = 8'b01000100; // **   **
         20'h00519: data = 8'b01010100; // ** * **
         20'h0051a: data = 8'b01011100; // ** ****
         20'h0051b: data = 8'b01111100; //  *****
         20'h0051c: data = 8'b00001100; //     **
         20'h0051d: data = 8'b00001100; //     ***
         20'h0051e: data = 8'b00000000; // 
         20'h0051f: data = 8'b00000000; // 
         //code x52   
         20'h00520: data = 8'b00000000; // 
         20'h00521: data = 8'b00000000; // 
         20'h00522: data = 8'b01111100; // ******
         20'h00523: data = 8'b00100110; //  **  **
         20'h00524: data = 8'b00100110; //  **  **
         20'h00525: data = 8'b00100110; //  **  **
         20'h00526: data = 8'b00111100; //  *****
         20'h00527: data = 8'b00100100; //  ** **
         20'h00528: data = 8'b00100100; //  **  **
         20'h00529: data = 8'b00100100; //  **  **
         20'h0052a: data = 8'b00100100; //  **  **
         20'h0052b: data = 8'b00100110; // ***  **
         20'h0052c: data = 8'b00000000; // 
         20'h0052d: data = 8'b00000000; // 
         20'h0052e: data = 8'b00000000; // 
         20'h0052f: data = 8'b00000000; // 
         //code x53   
         20'h00530: data = 8'b00000000; // 
         20'h00531: data = 8'b00000000; // 
         20'h00532: data = 8'b01111100; //  *****
         20'h00533: data = 8'b01000100; // **   **
         20'h00534: data = 8'b01000100; // **   **
         20'h00535: data = 8'b01100000; //  **
         20'h00536: data = 8'b00111000; //   ***
         20'h00537: data = 8'b00001100; //     **
         20'h00538: data = 8'b00000100; //      **
         20'h00539: data = 8'b01000100; // **   **
         20'h0053a: data = 8'b01000100; // **   **
         20'h0053b: data = 8'b01111100; //  *****
         20'h0053c: data = 8'b00000000; // 
         20'h0053d: data = 8'b00000000; // 
         20'h0053e: data = 8'b00000000; // 
         20'h0053f: data = 8'b00000000; // 
         //code x54   
         20'h00540: data = 8'b00000000; // 
         20'h00541: data = 8'b00000000; // 
         20'h00542: data = 8'b01111111; // ********
         20'h00543: data = 8'b01011011; // ** ** **
         20'h00544: data = 8'b00011001; // *  **  *
         20'h00545: data = 8'b00011000; //    **
         20'h00546: data = 8'b00011000; //    **
         20'h00547: data = 8'b00011000; //    **
         20'h00548: data = 8'b00011000; //    **
         20'h00549: data = 8'b00011000; //    **
         20'h0054a: data = 8'b00011000; //    **
         20'h0054b: data = 8'b00111100; //   ****
         20'h0054c: data = 8'b00000000; // 
         20'h0054d: data = 8'b00000000; // 
         20'h0054e: data = 8'b00000000; // 
         20'h0054f: data = 8'b00000000; // 
         //code x55   
         20'h00550: data = 8'b00000000; // 
         20'h00551: data = 8'b00000000; // 
         20'h00552: data = 8'b01000100; // **   **
         20'h00553: data = 8'b01000100; // **   **
         20'h00554: data = 8'b01000100; // **   **
         20'h00555: data = 8'b01000100; // **   **
         20'h00556: data = 8'b01000100; // **   **
         20'h00557: data = 8'b01000100; // **   **
         20'h00558: data = 8'b01000100; // **   **
         20'h00559: data = 8'b01000100; // **   **
         20'h0055a: data = 8'b01000100; // **   **
         20'h0055b: data = 8'b01111100; //  *****
         20'h0055c: data = 8'b00000000; // 
         20'h0055d: data = 8'b00000000; // 
         20'h0055e: data = 8'b00000000; // 
         20'h0055f: data = 8'b00000000; // 
         //code x56   
         20'h00560: data = 8'b00000000; // 
         20'h00561: data = 8'b00000000; // 
         20'h00562: data = 8'b01000010; // **    **
         20'h00563: data = 8'b01000010; // **    **
         20'h00564: data = 8'b01000010; // **    **
         20'h00565: data = 8'b01000010; // **    **
         20'h00566: data = 8'b01000010; // **    **
         20'h00567: data = 8'b01000010; // **    **
         20'h00568: data = 8'b01000010; // **    **
         20'h00569: data = 8'b01100100; //  **  **
         20'h0056a: data = 8'b00111100; //   ****
         20'h0056b: data = 8'b00011000; //    **
         20'h0056c: data = 8'b00000000; // 
         20'h0056d: data = 8'b00000000; // 
         20'h0056e: data = 8'b00000000; // 
         20'h0056f: data = 8'b00000000; // 
         //code x57   
         20'h00570: data = 8'b00000000; // 
         20'h00571: data = 8'b00000000; // 
         20'h00572: data = 8'b01000010; // **    **
         20'h00573: data = 8'b01000010; // **    **
         20'h00574: data = 8'b01000010; // **    **
         20'h00575: data = 8'b01000010; // **    **
         20'h00576: data = 8'b01000010; // **    **
         20'h00577: data = 8'b01011010; // ** ** **
         20'h00578: data = 8'b01011010; // ** ** **
         20'h00579: data = 8'b01111110; // ********
         20'h0057a: data = 8'b01100100; //  **  **
         20'h0057b: data = 8'b01100100; //  **  **
         20'h0057c: data = 8'b00000000; // 
         20'h0057d: data = 8'b00000000; // 
         20'h0057e: data = 8'b00000000; // 
         20'h0057f: data = 8'b00000000; // 
         //code x58   
         20'h00580: data = 8'b00000000; // 
         20'h00581: data = 8'b00000000; // 
         20'h00582: data = 8'b01000011; // **    **
         20'h00583: data = 8'b01000011; // **    **
         20'h00584: data = 8'b01100100; //  **  **
         20'h00585: data = 8'b00111100; //   ****
         20'h00586: data = 8'b00011000; //    **
         20'h00587: data = 8'b00011000; //    **
         20'h00588: data = 8'b00111100; //   ****
         20'h00589: data = 8'b01100100; //  **  **
         20'h0058a: data = 8'b01000011; // **    **
         20'h0058b: data = 8'b01000011; // **    **
         20'h0058c: data = 8'b00000000; // 
         20'h0058d: data = 8'b00000000; // 
         20'h0058e: data = 8'b00000000; // 
         20'h0058f: data = 8'b00000000; // 
         //code x59   
         20'h00590: data = 8'b00000000; // 
         20'h00591: data = 8'b00000000; // 
         20'h00592: data = 8'b01000011; // **    **
         20'h00593: data = 8'b01000011; // **    **
         20'h00594: data = 8'b01000011; // **    **
         20'h00595: data = 8'b01100100; //  **  **
         20'h00596: data = 8'b00111100; //   ****
         20'h00597: data = 8'b00011000; //    **
         20'h00598: data = 8'b00011000; //    **
         20'h00599: data = 8'b00011000; //    **
         20'h0059a: data = 8'b00011000; //    **
         20'h0059b: data = 8'b00111100; //   ****
         20'h0059c: data = 8'b00000000; // 
         20'h0059d: data = 8'b00000000; // 
         20'h0059e: data = 8'b00000000; // 
         20'h0059f: data = 8'b00000000; // 
         //code x5a   
         20'h005a0: data = 8'b00000000; // 
         20'h005a1: data = 8'b00000000; // 
         20'h005a2: data = 8'b01111111; // ********
         20'h005a3: data = 8'b01000011; // **    **
         20'h005a4: data = 8'b00000100; // *    **
         20'h005a5: data = 8'b00001100; //     **
         20'h005a6: data = 8'b00011000; //    **
         20'h005a7: data = 8'b00110000; //   **
         20'h005a8: data = 8'b01100000; //  **
         20'h005a9: data = 8'b01000001; // **     *
         20'h005aa: data = 8'b01000011; // **    **
         20'h005ab: data = 8'b01111111; // ********
         20'h005ac: data = 8'b00000000; // 
         20'h005ad: data = 8'b00000000; // 
         20'h005ae: data = 8'b00000000; // 
         20'h005af: data = 8'b00000000; // 
         //code x5b   
         20'h005b0: data = 8'b00000000; // 
         20'h005b1: data = 8'b00000000; // 
         20'h005b2: data = 8'b00111100; //   ****
         20'h005b3: data = 8'b00110000; //   **
         20'h005b4: data = 8'b00110000; //   **
         20'h005b5: data = 8'b00110000; //   **
         20'h005b6: data = 8'b00110000; //   **
         20'h005b7: data = 8'b00110000; //   **
         20'h005b8: data = 8'b00110000; //   **
         20'h005b9: data = 8'b00110000; //   **
         20'h005ba: data = 8'b00110000; //   **
         20'h005bb: data = 8'b00111100; //   ****
         20'h005bc: data = 8'b00000000; // 
         20'h005bd: data = 8'b00000000; // 
         20'h005be: data = 8'b00000000; // 
         20'h005bf: data = 8'b00000000; // 
         //code x5c   
         20'h005c0: data = 8'b00000000; // 
         20'h005c1: data = 8'b00000000; // 
         20'h005c2: data = 8'b00000000; // 
         20'h005c3: data = 8'b00000000; // *
         20'h005c4: data = 8'b01000000; // **
         20'h005c5: data = 8'b01100000; // ***
         20'h005c6: data = 8'b01110000; //  ***
         20'h005c7: data = 8'b00111000; //   ***
         20'h005c8: data = 8'b00011100; //    ***
         20'h005c9: data = 8'b00001100; //     ***
         20'h005ca: data = 8'b00000100; //      **
         20'h005cb: data = 8'b00000000; //       *
         20'h005cc: data = 8'b00000000; // 
         20'h005cd: data = 8'b00000000; // 
         20'h005ce: data = 8'b00000000; // 
         20'h005cf: data = 8'b00000000; // 
         //code x5d   
         20'h005d0: data = 8'b00000000; // 
         20'h005d1: data = 8'b00000000; // 
         20'h005d2: data = 8'b00111100; //   ****
         20'h005d3: data = 8'b00001100; //     **
         20'h005d4: data = 8'b00001100; //     **
         20'h005d5: data = 8'b00001100; //     **
         20'h005d6: data = 8'b00001100; //     **
         20'h005d7: data = 8'b00001100; //     **
         20'h005d8: data = 8'b00001100; //     **
         20'h005d9: data = 8'b00001100; //     **
         20'h005da: data = 8'b00001100; //     **
         20'h005db: data = 8'b00111100; //   ****
         20'h005dc: data = 8'b00000000; // 
         20'h005dd: data = 8'b00000000; // 
         20'h005de: data = 8'b00000000; // 
         20'h005df: data = 8'b00000000; // 
         //code x5e   
         20'h005e0: data = 8'b00010000; //    *
         20'h005e1: data = 8'b00111000; //   ***
         20'h005e2: data = 8'b01101100; //  ** **
         20'h005e3: data = 8'b01000100; // **   **
         20'h005e4: data = 8'b00000000; // 
         20'h005e5: data = 8'b00000000; // 
         20'h005e6: data = 8'b00000000; // 
         20'h005e7: data = 8'b00000000; // 
         20'h005e8: data = 8'b00000000; // 
         20'h005e9: data = 8'b00000000; // 
         20'h005ea: data = 8'b00000000; // 
         20'h005eb: data = 8'b00000000; // 
         20'h005ec: data = 8'b00000000; // 
         20'h005ed: data = 8'b00000000; // 
         20'h005ee: data = 8'b00000000; // 
         20'h005ef: data = 8'b00000000; // 
         //code x5f   
         20'h005f0: data = 8'b00000000; // 
         20'h005f1: data = 8'b00000000; // 
         20'h005f2: data = 8'b00000000; // 
         20'h005f3: data = 8'b00000000; // 
         20'h005f4: data = 8'b00000000; // 
         20'h005f5: data = 8'b00000000; // 
         20'h005f6: data = 8'b00000000; // 
         20'h005f7: data = 8'b00000000; // 
         20'h005f8: data = 8'b00000000; // 
         20'h005f9: data = 8'b00000000; // 
         20'h005fa: data = 8'b00000000; // 
         20'h005fb: data = 8'b00000000; // 
         20'h005fc: data = 8'b00000000; // 
         20'h005fd: data = 8'b01111111; // ********
         20'h005fe: data = 8'b00000000; // 
         20'h005ff: data = 8'b00000000; // 
         //code x60   
         20'h00600: data = 8'b00110000; //   **
         20'h00601: data = 8'b00110000; //   **
         20'h00602: data = 8'b00011000; //    **
         20'h00603: data = 8'b00000000; // 
         20'h00604: data = 8'b00000000; // 
         20'h00605: data = 8'b00000000; // 
         20'h00606: data = 8'b00000000; // 
         20'h00607: data = 8'b00000000; // 
         20'h00608: data = 8'b00000000; // 
         20'h00609: data = 8'b00000000; // 
         20'h0060a: data = 8'b00000000; // 
         20'h0060b: data = 8'b00000000; // 
         20'h0060c: data = 8'b00000000; // 
         20'h0060d: data = 8'b00000000; // 
         20'h0060e: data = 8'b00000000; // 
         20'h0060f: data = 8'b00000000; // 
         //code x61   
         20'h00610: data = 8'b00000000; // 
         20'h00611: data = 8'b00000000; // 
         20'h00612: data = 8'b00000000; // 
         20'h00613: data = 8'b00000000; // 
         20'h00614: data = 8'b00000000; // 
         20'h00615: data = 8'b01111000; //  ****
         20'h00616: data = 8'b00001100; //     **
         20'h00617: data = 8'b01111100; //  *****
         20'h00618: data = 8'b01001100; // **  **
         20'h00619: data = 8'b01001100; // **  **
         20'h0061a: data = 8'b01001100; // **  **
         20'h0061b: data = 8'b01110100; //  *** **
         20'h0061c: data = 8'b00000000; // 
         20'h0061d: data = 8'b00000000; // 
         20'h0061e: data = 8'b00000000; // 
         20'h0061f: data = 8'b00000000; // 
         //code x62   
         20'h00620: data = 8'b00000000; // 
         20'h00621: data = 8'b00000000; // 
         20'h00622: data = 8'b01100000; //  ***
         20'h00623: data = 8'b01100000; //   **
         20'h00624: data = 8'b01100000; //   **
         20'h00625: data = 8'b01111000; //   ****
         20'h00626: data = 8'b01101100; //   ** **
         20'h00627: data = 8'b01100100; //   **  **
         20'h00628: data = 8'b01100100; //   **  **
         20'h00629: data = 8'b01100100; //   **  **
         20'h0062a: data = 8'b01100100; //   **  **
         20'h0062b: data = 8'b01111100; //   *****
         20'h0062c: data = 8'b00000000; // 
         20'h0062d: data = 8'b00000000; // 
         20'h0062e: data = 8'b00000000; // 
         20'h0062f: data = 8'b00000000; // 
         //code x63   
         20'h00630: data = 8'b00000000; // 
         20'h00631: data = 8'b00000000; // 
         20'h00632: data = 8'b00000000; // 
         20'h00633: data = 8'b00000000; // 
         20'h00634: data = 8'b00000000; // 
         20'h00635: data = 8'b01111100; //  *****
         20'h00636: data = 8'b01000100; // **   **
         20'h00637: data = 8'b01000000; // **
         20'h00638: data = 8'b01000000; // **
         20'h00639: data = 8'b01000000; // **
         20'h0063a: data = 8'b01000100; // **   **
         20'h0063b: data = 8'b01111100; //  *****
         20'h0063c: data = 8'b00000000; // 
         20'h0063d: data = 8'b00000000; // 
         20'h0063e: data = 8'b00000000; // 
         20'h0063f: data = 8'b00000000; // 
         //code x64   
         20'h00640: data = 8'b00000000; // 
         20'h00641: data = 8'b00000000; // 
         20'h00642: data = 8'b00011100; //    ***
         20'h00643: data = 8'b00001100; //     **
         20'h00644: data = 8'b00001100; //     **
         20'h00645: data = 8'b00111100; //   ****
         20'h00646: data = 8'b01101100; //  ** **
         20'h00647: data = 8'b01001100; // **  **
         20'h00648: data = 8'b01001100; // **  **
         20'h00649: data = 8'b01001100; // **  **
         20'h0064a: data = 8'b01001100; // **  **
         20'h0064b: data = 8'b01110100; //  *** **
         20'h0064c: data = 8'b00000000; // 
         20'h0064d: data = 8'b00000000; // 
         20'h0064e: data = 8'b00000000; // 
         20'h0064f: data = 8'b00000000; // 
         //code x65   
         20'h00650: data = 8'b00000000; // 
         20'h00651: data = 8'b00000000; // 
         20'h00652: data = 8'b00000000; // 
         20'h00653: data = 8'b00000000; // 
         20'h00654: data = 8'b00000000; // 
         20'h00655: data = 8'b01111100; //  *****
         20'h00656: data = 8'b01000100; // **   **
         20'h00657: data = 8'b01111100; // *******
         20'h00658: data = 8'b01000000; // **
         20'h00659: data = 8'b01000000; // **
         20'h0065a: data = 8'b01000100; // **   **
         20'h0065b: data = 8'b01111100; //  *****
         20'h0065c: data = 8'b00000000; // 
         20'h0065d: data = 8'b00000000; // 
         20'h0065e: data = 8'b00000000; // 
         20'h0065f: data = 8'b00000000; // 
         //code x66   
         20'h00660: data = 8'b00000000; // 
         20'h00661: data = 8'b00000000; // 
         20'h00662: data = 8'b00111000; //   ***
         20'h00663: data = 8'b01101100; //  ** **
         20'h00664: data = 8'b01100100; //  **  *
         20'h00665: data = 8'b01100000; //  **
         20'h00666: data = 8'b01110000; // ****
         20'h00667: data = 8'b01100000; //  **
         20'h00668: data = 8'b01100000; //  **
         20'h00669: data = 8'b01100000; //  **
         20'h0066a: data = 8'b01100000; //  **
         20'h0066b: data = 8'b01110000; // ****
         20'h0066c: data = 8'b00000000; // 
         20'h0066d: data = 8'b00000000; // 
         20'h0066e: data = 8'b00000000; // 
         20'h0066f: data = 8'b00000000; // 
         //code x67   
         20'h00670: data = 8'b00000000; // 
         20'h00671: data = 8'b00000000; // 
         20'h00672: data = 8'b00000000; // 
         20'h00673: data = 8'b00000000; // 
         20'h00674: data = 8'b00000000; // 
         20'h00675: data = 8'b01110100; //  *** **
         20'h00676: data = 8'b01001100; // **  **
         20'h00677: data = 8'b01001100; // **  **
         20'h00678: data = 8'b01001100; // **  **
         20'h00679: data = 8'b01001100; // **  **
         20'h0067a: data = 8'b01001100; // **  **
         20'h0067b: data = 8'b01111100; //  *****
         20'h0067c: data = 8'b00001100; //     **
         20'h0067d: data = 8'b01001100; // **  **
         20'h0067e: data = 8'b01111000; //  ****
         20'h0067f: data = 8'b00000000; // 
         //code x68   
         20'h00680: data = 8'b00000000; // 
         20'h00681: data = 8'b00000000; // 
         20'h00682: data = 8'b01100000; // ***
         20'h00683: data = 8'b01100000; //  **
         20'h00684: data = 8'b01100000; //  **
         20'h00685: data = 8'b01101100; //  ** **
         20'h00686: data = 8'b01110100; //  *** **
         20'h00687: data = 8'b01100100; //  **  **
         20'h00688: data = 8'b01100100; //  **  **
         20'h00689: data = 8'b01100100; //  **  **
         20'h0068a: data = 8'b01100100; //  **  **
         20'h0068b: data = 8'b01100100; // ***  **
         20'h0068c: data = 8'b00000000; // 
         20'h0068d: data = 8'b00000000; // 
         20'h0068e: data = 8'b00000000; // 
         20'h0068f: data = 8'b00000000; // 
         //code x69   
         20'h00690: data = 8'b00000000; // 
         20'h00691: data = 8'b00000000; // 
         20'h00692: data = 8'b00011000; //    **
         20'h00693: data = 8'b00011000; //    **
         20'h00694: data = 8'b00000000; // 
         20'h00695: data = 8'b00111000; //   ***
         20'h00696: data = 8'b00011000; //    **
         20'h00697: data = 8'b00011000; //    **
         20'h00698: data = 8'b00011000; //    **
         20'h00699: data = 8'b00011000; //    **
         20'h0069a: data = 8'b00011000; //    **
         20'h0069b: data = 8'b00111100; //   ****
         20'h0069c: data = 8'b00000000; // 
         20'h0069d: data = 8'b00000000; // 
         20'h0069e: data = 8'b00000000; // 
         20'h0069f: data = 8'b00000000; // 
         //code x6a   
         20'h006a0: data = 8'b00000000; // 
         20'h006a1: data = 8'b00000000; // 
         20'h006a2: data = 8'b00000100; //      **
         20'h006a3: data = 8'b00000100; //      **
         20'h006a4: data = 8'b00000000; // 
         20'h006a5: data = 8'b00001100; //     ***
         20'h006a6: data = 8'b00000100; //      **
         20'h006a7: data = 8'b00000100; //      **
         20'h006a8: data = 8'b00000100; //      **
         20'h006a9: data = 8'b00000100; //      **
         20'h006aa: data = 8'b00000100; //      **
         20'h006ab: data = 8'b00000100; //      **
         20'h006ac: data = 8'b01100100; //  **  **
         20'h006ad: data = 8'b01100100; //  **  **
         20'h006ae: data = 8'b00111100; //   ****
         20'h006af: data = 8'b00000000; // 
         //code x6b   
         20'h006b0: data = 8'b00000000; // 
         20'h006b1: data = 8'b00000000; // 
         20'h006b2: data = 8'b01100000; // ***
         20'h006b3: data = 8'b01100000; //  **
         20'h006b4: data = 8'b01100000; //  **
         20'h006b5: data = 8'b01100100; //  **  **
         20'h006b6: data = 8'b01101100; //  ** **
         20'h006b7: data = 8'b01111000; //  ****
         20'h006b8: data = 8'b01111000; //  ****
         20'h006b9: data = 8'b01101100; //  ** **
         20'h006ba: data = 8'b01100100; //  **  **
         20'h006bb: data = 8'b01100100; // ***  **
         20'h006bc: data = 8'b00000000; // 
         20'h006bd: data = 8'b00000000; // 
         20'h006be: data = 8'b00000000; // 
         20'h006bf: data = 8'b00000000; // 
         //code x6c   
         20'h006c0: data = 8'b00000000; // 
         20'h006c1: data = 8'b00000000; // 
         20'h006c2: data = 8'b00111000; //   ***
         20'h006c3: data = 8'b00011000; //    **
         20'h006c4: data = 8'b00011000; //    **
         20'h006c5: data = 8'b00011000; //    **
         20'h006c6: data = 8'b00011000; //    **
         20'h006c7: data = 8'b00011000; //    **
         20'h006c8: data = 8'b00011000; //    **
         20'h006c9: data = 8'b00011000; //    **
         20'h006ca: data = 8'b00011000; //    **
         20'h006cb: data = 8'b00111100; //   ****
         20'h006cc: data = 8'b00000000; // 
         20'h006cd: data = 8'b00000000; // 
         20'h006ce: data = 8'b00000000; // 
         20'h006cf: data = 8'b00000000; // 
         //code x6d   
         20'h006d0: data = 8'b00000000; // 
         20'h006d1: data = 8'b00000000; // 
         20'h006d2: data = 8'b00000000; // 
         20'h006d3: data = 8'b00000000; // 
         20'h006d4: data = 8'b00000000; // 
         20'h006d5: data = 8'b01100100; // ***  **
         20'h006d6: data = 8'b01111111; // ********
         20'h006d7: data = 8'b01011011; // ** ** **
         20'h006d8: data = 8'b01011011; // ** ** **
         20'h006d9: data = 8'b01011011; // ** ** **
         20'h006da: data = 8'b01011011; // ** ** **
         20'h006db: data = 8'b01011011; // ** ** **
         20'h006dc: data = 8'b00000000; // 
         20'h006dd: data = 8'b00000000; // 
         20'h006de: data = 8'b00000000; // 
         20'h006df: data = 8'b00000000; // 
         //code x6e   
         20'h006e0: data = 8'b00000000; // 
         20'h006e1: data = 8'b00000000; // 
         20'h006e2: data = 8'b00000000; // 
         20'h006e3: data = 8'b00000000; // 
         20'h006e4: data = 8'b00000000; // 
         20'h006e5: data = 8'b01011100; // ** ***
         20'h006e6: data = 8'b01100100; //  **  **
         20'h006e7: data = 8'b01100100; //  **  **
         20'h006e8: data = 8'b01100100; //  **  **
         20'h006e9: data = 8'b01100100; //  **  **
         20'h006ea: data = 8'b01100100; //  **  **
         20'h006eb: data = 8'b01100100; //  **  **
         20'h006ec: data = 8'b00000000; // 
         20'h006ed: data = 8'b00000000; // 
         20'h006ee: data = 8'b00000000; // 
         20'h006ef: data = 8'b00000000; // 
         //code x6f   
         20'h006f0: data = 8'b00000000; // 
         20'h006f1: data = 8'b00000000; // 
         20'h006f2: data = 8'b00000000; // 
         20'h006f3: data = 8'b00000000; // 
         20'h006f4: data = 8'b00000000; // 
         20'h006f5: data = 8'b01111100; //  *****
         20'h006f6: data = 8'b01000100; // **   **
         20'h006f7: data = 8'b01000100; // **   **
         20'h006f8: data = 8'b01000100; // **   **
         20'h006f9: data = 8'b01000100; // **   **
         20'h006fa: data = 8'b01000100; // **   **
         20'h006fb: data = 8'b01111100; //  *****
         20'h006fc: data = 8'b00000000; // 
         20'h006fd: data = 8'b00000000; // 
         20'h006fe: data = 8'b00000000; // 
         20'h006ff: data = 8'b00000000; // 
         //code x70   
         20'h00700: data = 8'b00000000; // 
         20'h00701: data = 8'b00000000; // 
         20'h00702: data = 8'b00000000; // 
         20'h00703: data = 8'b00000000; // 
         20'h00704: data = 8'b00000000; // 
         20'h00705: data = 8'b01011100; // ** ***
         20'h00706: data = 8'b01100100; //  **  **
         20'h00707: data = 8'b01100100; //  **  **
         20'h00708: data = 8'b01100100; //  **  **
         20'h00709: data = 8'b01100100; //  **  **
         20'h0070a: data = 8'b01100100; //  **  **
         20'h0070b: data = 8'b01111100; //  *****
         20'h0070c: data = 8'b01100000; //  **
         20'h0070d: data = 8'b01100000; //  **
         20'h0070e: data = 8'b01110000; // ****
         20'h0070f: data = 8'b00000000; // 
         //code x71   
         20'h00710: data = 8'b00000000; // 
         20'h00711: data = 8'b00000000; // 
         20'h00712: data = 8'b00000000; // 
         20'h00713: data = 8'b00000000; // 
         20'h00714: data = 8'b00000000; // 
         20'h00715: data = 8'b01110100; //  *** **
         20'h00716: data = 8'b01001100; // **  **
         20'h00717: data = 8'b01001100; // **  **
         20'h00718: data = 8'b01001100; // **  **
         20'h00719: data = 8'b01001100; // **  **
         20'h0071a: data = 8'b01001100; // **  **
         20'h0071b: data = 8'b01111100; //  *****
         20'h0071c: data = 8'b00001100; //     **
         20'h0071d: data = 8'b00001100; //     **
         20'h0071e: data = 8'b00011100; //    ****
         20'h0071f: data = 8'b00000000; // 
         //code x72   
         20'h00720: data = 8'b00000000; // 
         20'h00721: data = 8'b00000000; // 
         20'h00722: data = 8'b00000000; // 
         20'h00723: data = 8'b00000000; // 
         20'h00724: data = 8'b00000000; // 
         20'h00725: data = 8'b01011100; // ** ***
         20'h00726: data = 8'b01110100; //  *** **
         20'h00727: data = 8'b01100100; //  **  **
         20'h00728: data = 8'b01100000; //  **
         20'h00729: data = 8'b01100000; //  **
         20'h0072a: data = 8'b01100000; //  **
         20'h0072b: data = 8'b01110000; // ****
         20'h0072c: data = 8'b00000000; // 
         20'h0072d: data = 8'b00000000; // 
         20'h0072e: data = 8'b00000000; // 
         20'h0072f: data = 8'b00000000; // 
         //code x73   
         20'h00730: data = 8'b00000000; // 
         20'h00731: data = 8'b00000000; // 
         20'h00732: data = 8'b00000000; // 
         20'h00733: data = 8'b00000000; // 
         20'h00734: data = 8'b00000000; // 
         20'h00735: data = 8'b01111100; //  *****
         20'h00736: data = 8'b01000100; // **   **
         20'h00737: data = 8'b01100000; //  **
         20'h00738: data = 8'b00111000; //   ***
         20'h00739: data = 8'b00001100; //     **
         20'h0073a: data = 8'b01000100; // **   **
         20'h0073b: data = 8'b01111100; //  *****
         20'h0073c: data = 8'b00000000; // 
         20'h0073d: data = 8'b00000000; // 
         20'h0073e: data = 8'b00000000; // 
         20'h0073f: data = 8'b00000000; // 
         //code x74   
         20'h00740: data = 8'b00000000; // 
         20'h00741: data = 8'b00000000; // 
         20'h00742: data = 8'b00010000; //    *
         20'h00743: data = 8'b00110000; //   **
         20'h00744: data = 8'b00110000; //   **
         20'h00745: data = 8'b01111100; // ******
         20'h00746: data = 8'b00110000; //   **
         20'h00747: data = 8'b00110000; //   **
         20'h00748: data = 8'b00110000; //   **
         20'h00749: data = 8'b00110000; //   **
         20'h0074a: data = 8'b00110100; //   ** **
         20'h0074b: data = 8'b00011100; //    ***
         20'h0074c: data = 8'b00000000; // 
         20'h0074d: data = 8'b00000000; // 
         20'h0074e: data = 8'b00000000; // 
         20'h0074f: data = 8'b00000000; // 
         //code x75   
         20'h00750: data = 8'b00000000; // 
         20'h00751: data = 8'b00000000; // 
         20'h00752: data = 8'b00000000; // 
         20'h00753: data = 8'b00000000; // 
         20'h00754: data = 8'b00000000; // 
         20'h00755: data = 8'b01001100; // **  **
         20'h00756: data = 8'b01001100; // **  **
         20'h00757: data = 8'b01001100; // **  **
         20'h00758: data = 8'b01001100; // **  **
         20'h00759: data = 8'b01001100; // **  **
         20'h0075a: data = 8'b01001100; // **  **
         20'h0075b: data = 8'b01110100; //  *** **
         20'h0075c: data = 8'b00000000; // 
         20'h0075d: data = 8'b00000000; // 
         20'h0075e: data = 8'b00000000; // 
         20'h0075f: data = 8'b00000000; // 
         //code x76   
         20'h00760: data = 8'b00000000; // 
         20'h00761: data = 8'b00000000; // 
         20'h00762: data = 8'b00000000; // 
         20'h00763: data = 8'b00000000; // 
         20'h00764: data = 8'b00000000; // 
         20'h00765: data = 8'b01000011; // **    **
         20'h00766: data = 8'b01000011; // **    **
         20'h00767: data = 8'b01000011; // **    **
         20'h00768: data = 8'b01000011; // **    **
         20'h00769: data = 8'b01100100; //  **  **
         20'h0076a: data = 8'b00111100; //   ****
         20'h0076b: data = 8'b00011000; //    **
         20'h0076c: data = 8'b00000000; // 
         20'h0076d: data = 8'b00000000; // 
         20'h0076e: data = 8'b00000000; // 
         20'h0076f: data = 8'b00000000; // 
         //code x77   
         20'h00770: data = 8'b00000000; // 
         20'h00771: data = 8'b00000000; // 
         20'h00772: data = 8'b00000000; // 
         20'h00773: data = 8'b00000000; // 
         20'h00774: data = 8'b00000000; // 
         20'h00775: data = 8'b01000011; // **    **
         20'h00776: data = 8'b01000011; // **    **
         20'h00777: data = 8'b01000011; // **    **
         20'h00778: data = 8'b01011011; // ** ** **
         20'h00779: data = 8'b01011011; // ** ** **
         20'h0077a: data = 8'b01111111; // ********
         20'h0077b: data = 8'b01100100; //  **  **
         20'h0077c: data = 8'b00000000; // 
         20'h0077d: data = 8'b00000000; // 
         20'h0077e: data = 8'b00000000; // 
         20'h0077f: data = 8'b00000000; // 
         //code x78   
         20'h00780: data = 8'b00000000; // 
         20'h00781: data = 8'b00000000; // 
         20'h00782: data = 8'b00000000; // 
         20'h00783: data = 8'b00000000; // 
         20'h00784: data = 8'b00000000; // 
         20'h00785: data = 8'b01000011; // **    **
         20'h00786: data = 8'b01100100; //  **  **
         20'h00787: data = 8'b00111100; //   ****
         20'h00788: data = 8'b00011000; //    **
         20'h00789: data = 8'b00111100; //   ****
         20'h0078a: data = 8'b01100100; //  **  **
         20'h0078b: data = 8'b01000011; // **    **
         20'h0078c: data = 8'b00000000; // 
         20'h0078d: data = 8'b00000000; // 
         20'h0078e: data = 8'b00000000; // 
         20'h0078f: data = 8'b00000000; // 
         //code x79   
         20'h00790: data = 8'b00000000; // 
         20'h00791: data = 8'b00000000; // 
         20'h00792: data = 8'b00000000; // 
         20'h00793: data = 8'b00000000; // 
         20'h00794: data = 8'b00000000; // 
         20'h00795: data = 8'b01000100; // **   **
         20'h00796: data = 8'b01000100; // **   **
         20'h00797: data = 8'b01000100; // **   **
         20'h00798: data = 8'b01000100; // **   **
         20'h00799: data = 8'b01000100; // **   **
         20'h0079a: data = 8'b01000100; // **   **
         20'h0079b: data = 8'b01111100; //  ******
         20'h0079c: data = 8'b00000100; //      **
         20'h0079d: data = 8'b00001100; //     **
         20'h0079e: data = 8'b01111000; // *****
         20'h0079f: data = 8'b00000000; // 
         //code x7a   
         20'h007a0: data = 8'b00000000; // 
         20'h007a1: data = 8'b00000000; // 
         20'h007a2: data = 8'b00000000; // 
         20'h007a3: data = 8'b00000000; // 
         20'h007a4: data = 8'b00000000; // 
         20'h007a5: data = 8'b01111100; // *******
         20'h007a6: data = 8'b01001100; // **  **
         20'h007a7: data = 8'b00011000; //    **
         20'h007a8: data = 8'b00110000; //   **
         20'h007a9: data = 8'b01100000; //  **
         20'h007aa: data = 8'b01000100; // **   **
         20'h007ab: data = 8'b01111100; // *******
         20'h007ac: data = 8'b00000000; // 
         20'h007ad: data = 8'b00000000; // 
         20'h007ae: data = 8'b00000000; // 
         20'h007af: data = 8'b00000000; // 
         //code x7b   
         20'h007b0: data = 8'b00000000; // 
         20'h007b1: data = 8'b00000000; // 
         20'h007b2: data = 8'b00001100; //     ***
         20'h007b3: data = 8'b00011000; //    **
         20'h007b4: data = 8'b00011000; //    **
         20'h007b5: data = 8'b00011000; //    **
         20'h007b6: data = 8'b01110000; //  ***
         20'h007b7: data = 8'b00011000; //    **
         20'h007b8: data = 8'b00011000; //    **
         20'h007b9: data = 8'b00011000; //    **
         20'h007ba: data = 8'b00011000; //    **
         20'h007bb: data = 8'b00001100; //     ***
         20'h007bc: data = 8'b00000000; // 
         20'h007bd: data = 8'b00000000; // 
         20'h007be: data = 8'b00000000; // 
         20'h007bf: data = 8'b00000000; // 
         //code x7c   
         20'h007c0: data = 8'b00000000; // 
         20'h007c1: data = 8'b00000000; // 
         20'h007c2: data = 8'b00010000; //    **
         20'h007c3: data = 8'b00010000; //    **
         20'h007c4: data = 8'b00010000; //    **
         20'h007c5: data = 8'b00010000; //    **
         20'h007c6: data = 8'b00010000; // 
         20'h007c7: data = 8'b00010000; //    **
         20'h007c8: data = 8'b00010000; //    **
         20'h007c9: data = 8'b00010000; //    **
         20'h007ca: data = 8'b00010000; //    **
         20'h007cb: data = 8'b00010000; //    **
         20'h007cc: data = 8'b00000000; // 
         20'h007cd: data = 8'b00000000; // 
         20'h007ce: data = 8'b00000000; // 
         20'h007cf: data = 8'b00000000; // 
         //code x7d   
         20'h007d0: data = 8'b00000000; // 
         20'h007d1: data = 8'b00000000; // 
         20'h007d2: data = 8'b01110000; //  ***
         20'h007d3: data = 8'b00011000; //    **
         20'h007d4: data = 8'b00011000; //    **
         20'h007d5: data = 8'b00011000; //    **
         20'h007d6: data = 8'b00001100; //     ***
         20'h007d7: data = 8'b00011000; //    **
         20'h007d8: data = 8'b00011000; //    **
         20'h007d9: data = 8'b00011000; //    **
         20'h007da: data = 8'b00011000; //    **
         20'h007db: data = 8'b01110000; //  ***
         20'h007dc: data = 8'b00000000; // 
         20'h007dd: data = 8'b00000000; // 
         20'h007de: data = 8'b00000000; // 
         20'h007df: data = 8'b00000000; // 
         //code x7e   
         20'h007e0: data = 8'b00000000; // 
         20'h007e1: data = 8'b00000000; // 
         20'h007e2: data = 8'b01110100; //  *** **
         20'h007e3: data = 8'b01011100; // ** ***
         20'h007e4: data = 8'b00000000; // 
         20'h007e5: data = 8'b00000000; // 
         20'h007e6: data = 8'b00000000; // 
         20'h007e7: data = 8'b00000000; // 
         20'h007e8: data = 8'b00000000; // 
         20'h007e9: data = 8'b00000000; // 
         20'h007ea: data = 8'b00000000; // 
         20'h007eb: data = 8'b00000000; // 
         20'h007ec: data = 8'b00000000; // 
         20'h007ed: data = 8'b00000000; // 
         20'h007ee: data = 8'b00000000; // 
         20'h007ef: data = 8'b00000000; // 
         //code x7f   
         20'h007f0: data = 8'b00000000; // 
         20'h007f1: data = 8'b00000000; // 
         20'h007f2: data = 8'b00000000; // 
         20'h007f3: data = 8'b00000000; // 
         20'h007f4: data = 8'b00010000; //    *
         20'h007f5: data = 8'b00111000; //   ***
         20'h007f6: data = 8'b01101100; //  ** **
         20'h007f7: data = 8'b01000100; // **   **
         20'h007f8: data = 8'b01000100; // **   **
         20'h007f9: data = 8'b01000100; // **   **
         20'h007fa: data = 8'b01111100; // *******
         20'h007fb: data = 8'b00000000; // 
         20'h007fc: data = 8'b00000000; // 
         20'h007fd: data = 8'b00000000; // 
         20'h007fe: data = 8'b00000000; // 
         20'h007ff: data = 8'b00000000; //*/ 	 
   endcase
   
   always @(SELEC_PX,data[15],data[14],data[13],data[12],data[11],data[10],
   data[9],data[8], data[7], data[6], data[5], data[4], data[3], data[2], data[1], data[0])
      case (SELEC_PX)
      
         4'b0000: bit_fuente2 <= data[15];
         4'b0001: bit_fuente2 <= data[14]; 
         4'b0010: bit_fuente2 <= data[13];
         4'b0011: bit_fuente2 <= data[12];
         4'b0100: bit_fuente2 <= data[11];
         4'b0101: bit_fuente2 <= data[10];
         4'b0110: bit_fuente2 <= data[9];
         4'b0111: bit_fuente2 <= data[8];
	     4'b1000: bit_fuente2 <= data[7];
	     4'b1001: bit_fuente2 <= data[6];
	     4'b1010: bit_fuente2 <= data[5];
         4'b1011: bit_fuente2 <= data[4];
         4'b1100: bit_fuente2 <= data[3];
         4'b1101: bit_fuente2 <= data[2];
         4'b1110: bit_fuente2 <= data[1];
         4'b1111: bit_fuente2 <= data[0];
         default: bit_fuente2 <= 1'b0;
      endcase
   	     
   	     assign BIT_FUENTE2 = bit_fuente2;

endmodule      
	       